library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"ccfcc287",
    12 => x"86c0c84e",
    13 => x"49ccfcc2",
    14 => x"48ece4c2",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087c8e9",
    19 => x"1e87fc98",
    20 => x"1e731e72",
    21 => x"02114812",
    22 => x"c34b87ca",
    23 => x"739b98df",
    24 => x"87f00288",
    25 => x"4a264b26",
    26 => x"731e4f26",
    27 => x"c11e721e",
    28 => x"87ca048b",
    29 => x"02114812",
    30 => x"028887c4",
    31 => x"4a2687f1",
    32 => x"4f264b26",
    33 => x"731e741e",
    34 => x"c11e721e",
    35 => x"87d0048b",
    36 => x"02114812",
    37 => x"c34c87ca",
    38 => x"749c98df",
    39 => x"87eb0288",
    40 => x"4b264a26",
    41 => x"4f264c26",
    42 => x"8148731e",
    43 => x"c502a973",
    44 => x"05531287",
    45 => x"4f2687f6",
    46 => x"721e731e",
    47 => x"e7c0029a",
    48 => x"c148c087",
    49 => x"06a9724b",
    50 => x"827287d1",
    51 => x"7387c906",
    52 => x"01a97283",
    53 => x"87c387f4",
    54 => x"723ab2c1",
    55 => x"738903a9",
    56 => x"2ac10780",
    57 => x"87f3052b",
    58 => x"4f264b26",
    59 => x"c41e751e",
    60 => x"a1b7714d",
    61 => x"c1b9ff04",
    62 => x"07bdc381",
    63 => x"04a2b772",
    64 => x"82c1baff",
    65 => x"fe07bdc1",
    66 => x"2dc187ee",
    67 => x"c1b8ff04",
    68 => x"042d0780",
    69 => x"81c1b9ff",
    70 => x"264d2607",
    71 => x"4a711e4f",
    72 => x"484966c4",
    73 => x"a6c888c1",
    74 => x"02997158",
    75 => x"481287d4",
    76 => x"7808d4ff",
    77 => x"484966c4",
    78 => x"a6c888c1",
    79 => x"05997158",
    80 => x"4f2687ec",
    81 => x"c44a711e",
    82 => x"c1484966",
    83 => x"58a6c888",
    84 => x"d6029971",
    85 => x"48d4ff87",
    86 => x"6878ffc3",
    87 => x"4966c452",
    88 => x"c888c148",
    89 => x"997158a6",
    90 => x"2687ea05",
    91 => x"1e731e4f",
    92 => x"c34bd4ff",
    93 => x"4a6b7bff",
    94 => x"6b7bffc3",
    95 => x"7232c849",
    96 => x"7bffc3b1",
    97 => x"31c84a6b",
    98 => x"ffc3b271",
    99 => x"c8496b7b",
   100 => x"71b17232",
   101 => x"2687c448",
   102 => x"264c264d",
   103 => x"0e4f264b",
   104 => x"5d5c5b5e",
   105 => x"ff4a710e",
   106 => x"49724cd4",
   107 => x"7199ffc3",
   108 => x"ece4c27c",
   109 => x"87c805bf",
   110 => x"c94866d0",
   111 => x"58a6d430",
   112 => x"d84966d0",
   113 => x"99ffc329",
   114 => x"66d07c71",
   115 => x"c329d049",
   116 => x"7c7199ff",
   117 => x"c84966d0",
   118 => x"99ffc329",
   119 => x"66d07c71",
   120 => x"99ffc349",
   121 => x"49727c71",
   122 => x"ffc329d0",
   123 => x"6c7c7199",
   124 => x"fff0c94b",
   125 => x"abffc34d",
   126 => x"c387d005",
   127 => x"4b6c7cff",
   128 => x"c6028dc1",
   129 => x"abffc387",
   130 => x"7387f002",
   131 => x"87c7fe48",
   132 => x"ff49c01e",
   133 => x"ffc348d4",
   134 => x"c381c178",
   135 => x"04a9b7c8",
   136 => x"4f2687f1",
   137 => x"e71e731e",
   138 => x"dff8c487",
   139 => x"c01ec04b",
   140 => x"f7c1f0ff",
   141 => x"87e7fd49",
   142 => x"a8c186c4",
   143 => x"87eac005",
   144 => x"c348d4ff",
   145 => x"c0c178ff",
   146 => x"c0c0c0c0",
   147 => x"f0e1c01e",
   148 => x"fd49e9c1",
   149 => x"86c487c9",
   150 => x"ca059870",
   151 => x"48d4ff87",
   152 => x"c178ffc3",
   153 => x"fe87cb48",
   154 => x"8bc187e6",
   155 => x"87fdfe05",
   156 => x"e6fc48c0",
   157 => x"1e731e87",
   158 => x"c348d4ff",
   159 => x"4bd378ff",
   160 => x"ffc01ec0",
   161 => x"49c1c1f0",
   162 => x"c487d4fc",
   163 => x"05987086",
   164 => x"d4ff87ca",
   165 => x"78ffc348",
   166 => x"87cb48c1",
   167 => x"c187f1fd",
   168 => x"dbff058b",
   169 => x"fb48c087",
   170 => x"5e0e87f1",
   171 => x"ff0e5c5b",
   172 => x"dbfd4cd4",
   173 => x"1eeac687",
   174 => x"c1f0e1c0",
   175 => x"defb49c8",
   176 => x"c186c487",
   177 => x"87c802a8",
   178 => x"c087eafe",
   179 => x"87e2c148",
   180 => x"7087dafa",
   181 => x"ffffcf49",
   182 => x"a9eac699",
   183 => x"fe87c802",
   184 => x"48c087d3",
   185 => x"c387cbc1",
   186 => x"f1c07cff",
   187 => x"87f4fc4b",
   188 => x"c0029870",
   189 => x"1ec087eb",
   190 => x"c1f0ffc0",
   191 => x"defa49fa",
   192 => x"7086c487",
   193 => x"87d90598",
   194 => x"6c7cffc3",
   195 => x"7cffc349",
   196 => x"c17c7c7c",
   197 => x"c40299c0",
   198 => x"d548c187",
   199 => x"d148c087",
   200 => x"05abc287",
   201 => x"48c087c4",
   202 => x"8bc187c8",
   203 => x"87fdfe05",
   204 => x"e4f948c0",
   205 => x"1e731e87",
   206 => x"48ece4c2",
   207 => x"4bc778c1",
   208 => x"c248d0ff",
   209 => x"87c8fb78",
   210 => x"c348d0ff",
   211 => x"c01ec078",
   212 => x"c0c1d0e5",
   213 => x"87c7f949",
   214 => x"a8c186c4",
   215 => x"4b87c105",
   216 => x"c505abc2",
   217 => x"c048c087",
   218 => x"8bc187f9",
   219 => x"87d0ff05",
   220 => x"c287f7fc",
   221 => x"7058f0e4",
   222 => x"87cd0598",
   223 => x"ffc01ec1",
   224 => x"49d0c1f0",
   225 => x"c487d8f8",
   226 => x"48d4ff86",
   227 => x"c478ffc3",
   228 => x"e4c287de",
   229 => x"d0ff58f4",
   230 => x"ff78c248",
   231 => x"ffc348d4",
   232 => x"f748c178",
   233 => x"5e0e87f5",
   234 => x"0e5d5c5b",
   235 => x"ffc34a71",
   236 => x"4cd4ff4d",
   237 => x"d0ff7c75",
   238 => x"78c3c448",
   239 => x"1e727c75",
   240 => x"c1f0ffc0",
   241 => x"d6f749d8",
   242 => x"7086c487",
   243 => x"87c50298",
   244 => x"f0c048c1",
   245 => x"c37c7587",
   246 => x"c0c87cfe",
   247 => x"4966d41e",
   248 => x"c487faf4",
   249 => x"757c7586",
   250 => x"d87c757c",
   251 => x"754be0da",
   252 => x"99496c7c",
   253 => x"c187c505",
   254 => x"87f3058b",
   255 => x"d0ff7c75",
   256 => x"c078c248",
   257 => x"87cff648",
   258 => x"5c5b5e0e",
   259 => x"4b710e5d",
   260 => x"eec54cc0",
   261 => x"ff4adfcd",
   262 => x"ffc348d4",
   263 => x"c3496878",
   264 => x"c005a9fe",
   265 => x"4d7087fd",
   266 => x"cc029b73",
   267 => x"1e66d087",
   268 => x"cff44973",
   269 => x"d686c487",
   270 => x"48d0ff87",
   271 => x"c378d1c4",
   272 => x"66d07dff",
   273 => x"d488c148",
   274 => x"987058a6",
   275 => x"ff87f005",
   276 => x"ffc348d4",
   277 => x"9b737878",
   278 => x"ff87c505",
   279 => x"78d048d0",
   280 => x"c14c4ac1",
   281 => x"eefe058a",
   282 => x"f4487487",
   283 => x"731e87e9",
   284 => x"c04a711e",
   285 => x"48d4ff4b",
   286 => x"ff78ffc3",
   287 => x"c3c448d0",
   288 => x"48d4ff78",
   289 => x"7278ffc3",
   290 => x"f0ffc01e",
   291 => x"f449d1c1",
   292 => x"86c487cd",
   293 => x"d2059870",
   294 => x"1ec0c887",
   295 => x"fd4966cc",
   296 => x"86c487e6",
   297 => x"d0ff4b70",
   298 => x"7378c248",
   299 => x"87ebf348",
   300 => x"5c5b5e0e",
   301 => x"1ec00e5d",
   302 => x"c1f0ffc0",
   303 => x"def349c9",
   304 => x"c21ed287",
   305 => x"fc49f4e4",
   306 => x"86c887fe",
   307 => x"84c14cc0",
   308 => x"04acb7d2",
   309 => x"e4c287f8",
   310 => x"49bf97f4",
   311 => x"c199c0c3",
   312 => x"c005a9c0",
   313 => x"e4c287e7",
   314 => x"49bf97fb",
   315 => x"e4c231d0",
   316 => x"4abf97fc",
   317 => x"b17232c8",
   318 => x"97fde4c2",
   319 => x"71b14abf",
   320 => x"ffffcf4c",
   321 => x"84c19cff",
   322 => x"e7c134ca",
   323 => x"fde4c287",
   324 => x"c149bf97",
   325 => x"c299c631",
   326 => x"bf97fee4",
   327 => x"2ab7c74a",
   328 => x"e4c2b172",
   329 => x"4abf97f9",
   330 => x"c29dcf4d",
   331 => x"bf97fae4",
   332 => x"ca9ac34a",
   333 => x"fbe4c232",
   334 => x"c24bbf97",
   335 => x"c2b27333",
   336 => x"bf97fce4",
   337 => x"9bc0c34b",
   338 => x"732bb7c6",
   339 => x"c181c2b2",
   340 => x"70307148",
   341 => x"7548c149",
   342 => x"724d7030",
   343 => x"7184c14c",
   344 => x"b7c0c894",
   345 => x"87cc06ad",
   346 => x"2db734c1",
   347 => x"adb7c0c8",
   348 => x"87f4ff01",
   349 => x"def04874",
   350 => x"5b5e0e87",
   351 => x"f80e5d5c",
   352 => x"daedc286",
   353 => x"c278c048",
   354 => x"c01ed2e5",
   355 => x"87defb49",
   356 => x"987086c4",
   357 => x"c087c505",
   358 => x"87cec948",
   359 => x"7ec14dc0",
   360 => x"bfc5fac0",
   361 => x"c8e6c249",
   362 => x"4bc8714a",
   363 => x"7087fbea",
   364 => x"87c20598",
   365 => x"fac07ec0",
   366 => x"c249bfc1",
   367 => x"714ae4e6",
   368 => x"e5ea4bc8",
   369 => x"05987087",
   370 => x"7ec087c2",
   371 => x"fdc0026e",
   372 => x"d8ecc287",
   373 => x"edc24dbf",
   374 => x"7ebf9fd0",
   375 => x"ead6c548",
   376 => x"87c705a8",
   377 => x"bfd8ecc2",
   378 => x"6e87ce4d",
   379 => x"d5e9ca48",
   380 => x"87c502a8",
   381 => x"f1c748c0",
   382 => x"d2e5c287",
   383 => x"f949751e",
   384 => x"86c487ec",
   385 => x"c5059870",
   386 => x"c748c087",
   387 => x"fac087dc",
   388 => x"c249bfc1",
   389 => x"714ae4e6",
   390 => x"cde94bc8",
   391 => x"05987087",
   392 => x"edc287c8",
   393 => x"78c148da",
   394 => x"fac087da",
   395 => x"c249bfc5",
   396 => x"714ac8e6",
   397 => x"f1e84bc8",
   398 => x"02987087",
   399 => x"c087c5c0",
   400 => x"87e6c648",
   401 => x"97d0edc2",
   402 => x"d5c149bf",
   403 => x"cdc005a9",
   404 => x"d1edc287",
   405 => x"c249bf97",
   406 => x"c002a9ea",
   407 => x"48c087c5",
   408 => x"c287c7c6",
   409 => x"bf97d2e5",
   410 => x"e9c3487e",
   411 => x"cec002a8",
   412 => x"c3486e87",
   413 => x"c002a8eb",
   414 => x"48c087c5",
   415 => x"c287ebc5",
   416 => x"bf97dde5",
   417 => x"c0059949",
   418 => x"e5c287cc",
   419 => x"49bf97de",
   420 => x"c002a9c2",
   421 => x"48c087c5",
   422 => x"c287cfc5",
   423 => x"bf97dfe5",
   424 => x"d6edc248",
   425 => x"484c7058",
   426 => x"edc288c1",
   427 => x"e5c258da",
   428 => x"49bf97e0",
   429 => x"e5c28175",
   430 => x"4abf97e1",
   431 => x"a17232c8",
   432 => x"e7f1c27e",
   433 => x"c2786e48",
   434 => x"bf97e2e5",
   435 => x"58a6c848",
   436 => x"bfdaedc2",
   437 => x"87d4c202",
   438 => x"bfc1fac0",
   439 => x"e4e6c249",
   440 => x"4bc8714a",
   441 => x"7087c3e6",
   442 => x"c5c00298",
   443 => x"c348c087",
   444 => x"edc287f8",
   445 => x"c24cbfd2",
   446 => x"c25cfbf1",
   447 => x"bf97f7e5",
   448 => x"c231c849",
   449 => x"bf97f6e5",
   450 => x"c249a14a",
   451 => x"bf97f8e5",
   452 => x"7232d04a",
   453 => x"e5c249a1",
   454 => x"4abf97f9",
   455 => x"a17232d8",
   456 => x"9166c449",
   457 => x"bfe7f1c2",
   458 => x"eff1c281",
   459 => x"ffe5c259",
   460 => x"c84abf97",
   461 => x"fee5c232",
   462 => x"a24bbf97",
   463 => x"c0e6c24a",
   464 => x"d04bbf97",
   465 => x"4aa27333",
   466 => x"97c1e6c2",
   467 => x"9bcf4bbf",
   468 => x"a27333d8",
   469 => x"f3f1c24a",
   470 => x"eff1c25a",
   471 => x"8ac24abf",
   472 => x"f1c29274",
   473 => x"a17248f3",
   474 => x"87cac178",
   475 => x"97e4e5c2",
   476 => x"31c849bf",
   477 => x"97e3e5c2",
   478 => x"49a14abf",
   479 => x"59e2edc2",
   480 => x"bfdeedc2",
   481 => x"c731c549",
   482 => x"29c981ff",
   483 => x"59fbf1c2",
   484 => x"97e9e5c2",
   485 => x"32c84abf",
   486 => x"97e8e5c2",
   487 => x"4aa24bbf",
   488 => x"6e9266c4",
   489 => x"f7f1c282",
   490 => x"eff1c25a",
   491 => x"c278c048",
   492 => x"7248ebf1",
   493 => x"f1c278a1",
   494 => x"f1c248fb",
   495 => x"c278bfef",
   496 => x"c248fff1",
   497 => x"78bff3f1",
   498 => x"bfdaedc2",
   499 => x"87c9c002",
   500 => x"30c44874",
   501 => x"c9c07e70",
   502 => x"f7f1c287",
   503 => x"30c448bf",
   504 => x"edc27e70",
   505 => x"786e48de",
   506 => x"8ef848c1",
   507 => x"4c264d26",
   508 => x"4f264b26",
   509 => x"5c5b5e0e",
   510 => x"4a710e5d",
   511 => x"bfdaedc2",
   512 => x"7287cb02",
   513 => x"722bc74b",
   514 => x"9cffc14c",
   515 => x"4b7287c9",
   516 => x"4c722bc8",
   517 => x"c29cffc3",
   518 => x"83bfe7f1",
   519 => x"bffdf9c0",
   520 => x"87d902ab",
   521 => x"5bc1fac0",
   522 => x"1ed2e5c2",
   523 => x"fdf04973",
   524 => x"7086c487",
   525 => x"87c50598",
   526 => x"e6c048c0",
   527 => x"daedc287",
   528 => x"87d202bf",
   529 => x"91c44974",
   530 => x"81d2e5c2",
   531 => x"ffcf4d69",
   532 => x"9dffffff",
   533 => x"497487cb",
   534 => x"e5c291c2",
   535 => x"699f81d2",
   536 => x"fe48754d",
   537 => x"5e0e87c6",
   538 => x"0e5d5c5b",
   539 => x"4c7186f4",
   540 => x"87c5059c",
   541 => x"f5c348c0",
   542 => x"7ea4c887",
   543 => x"78c0486e",
   544 => x"c70266dc",
   545 => x"9766dc87",
   546 => x"87c505bf",
   547 => x"ddc348c0",
   548 => x"c11ec087",
   549 => x"87c9d049",
   550 => x"a6c886c4",
   551 => x"0266c458",
   552 => x"c287ffc0",
   553 => x"dc4ae2ed",
   554 => x"deff4966",
   555 => x"987087e1",
   556 => x"87eec002",
   557 => x"dc4a66c4",
   558 => x"4bcb4966",
   559 => x"87c4dfff",
   560 => x"dd029870",
   561 => x"c81ec087",
   562 => x"87c40266",
   563 => x"87c24dc0",
   564 => x"49754dc1",
   565 => x"c487cacf",
   566 => x"58a6c886",
   567 => x"ff0566c4",
   568 => x"66c487c1",
   569 => x"87c4c202",
   570 => x"6e81dc49",
   571 => x"c4786948",
   572 => x"81da4966",
   573 => x"9f4da4c4",
   574 => x"edc27d69",
   575 => x"d502bfda",
   576 => x"4966c487",
   577 => x"699f81d4",
   578 => x"ffffc049",
   579 => x"d0487199",
   580 => x"58a6cc30",
   581 => x"a6c887c5",
   582 => x"c878c048",
   583 => x"6d484966",
   584 => x"c07d7080",
   585 => x"49a4cc7c",
   586 => x"a4d0796d",
   587 => x"c479c049",
   588 => x"78c048a6",
   589 => x"c44aa4d4",
   590 => x"91c84966",
   591 => x"c049a172",
   592 => x"c4796d41",
   593 => x"80c14866",
   594 => x"c658a6c8",
   595 => x"ff04a8b7",
   596 => x"bf6e87e2",
   597 => x"722ac94a",
   598 => x"4af0c049",
   599 => x"87d8ddff",
   600 => x"c4c14a70",
   601 => x"797249a4",
   602 => x"87c248c1",
   603 => x"8ef448c0",
   604 => x"0e87f9f9",
   605 => x"5d5c5b5e",
   606 => x"9c4c710e",
   607 => x"87cac102",
   608 => x"6949a4c8",
   609 => x"87c2c102",
   610 => x"6c4a66d0",
   611 => x"a6d48249",
   612 => x"4d66d05a",
   613 => x"d6edc2b9",
   614 => x"baff4abf",
   615 => x"99719972",
   616 => x"87e4c002",
   617 => x"6b4ba4c4",
   618 => x"87c8f949",
   619 => x"edc27b70",
   620 => x"6c49bfd2",
   621 => x"757c7181",
   622 => x"d6edc2b9",
   623 => x"baff4abf",
   624 => x"99719972",
   625 => x"87dcff05",
   626 => x"dff87c75",
   627 => x"1e731e87",
   628 => x"029b4b71",
   629 => x"a3c887c7",
   630 => x"c5056949",
   631 => x"c048c087",
   632 => x"f1c287f7",
   633 => x"c44abfeb",
   634 => x"496949a3",
   635 => x"edc289c2",
   636 => x"7191bfd2",
   637 => x"edc24aa2",
   638 => x"6b49bfd6",
   639 => x"4aa27199",
   640 => x"5ac1fac0",
   641 => x"721e66c8",
   642 => x"87e2e949",
   643 => x"987086c4",
   644 => x"c087c405",
   645 => x"c187c248",
   646 => x"87d4f748",
   647 => x"711e731e",
   648 => x"c7029b4b",
   649 => x"49a3c887",
   650 => x"87c50569",
   651 => x"f7c048c0",
   652 => x"ebf1c287",
   653 => x"a3c44abf",
   654 => x"c2496949",
   655 => x"d2edc289",
   656 => x"a27191bf",
   657 => x"d6edc24a",
   658 => x"996b49bf",
   659 => x"c04aa271",
   660 => x"c85ac1fa",
   661 => x"49721e66",
   662 => x"c487cbe5",
   663 => x"05987086",
   664 => x"48c087c4",
   665 => x"48c187c2",
   666 => x"0e87c5f6",
   667 => x"5d5c5b5e",
   668 => x"7186f80e",
   669 => x"c47eff4c",
   670 => x"ffc148a6",
   671 => x"ffffffff",
   672 => x"d44bc078",
   673 => x"49734aa4",
   674 => x"a17291c8",
   675 => x"4866d849",
   676 => x"49708869",
   677 => x"adb7c04d",
   678 => x"c487cc04",
   679 => x"03adb766",
   680 => x"7e7387c5",
   681 => x"c15da6c8",
   682 => x"abb7c683",
   683 => x"87d3ff04",
   684 => x"8ef8486e",
   685 => x"0e87f5f4",
   686 => x"5d5c5b5e",
   687 => x"7186f00e",
   688 => x"48a6c47e",
   689 => x"ffffffc1",
   690 => x"c478ffff",
   691 => x"c078ff80",
   692 => x"6e4cc04d",
   693 => x"7483d44b",
   694 => x"7392c84a",
   695 => x"49754aa2",
   696 => x"a17391c8",
   697 => x"69486a49",
   698 => x"d0497088",
   699 => x"ad7459a6",
   700 => x"cc87cf02",
   701 => x"66c44966",
   702 => x"87c603a9",
   703 => x"c85ca6cc",
   704 => x"84c159a6",
   705 => x"04acb7c6",
   706 => x"c187c8ff",
   707 => x"adb7c685",
   708 => x"87fdfe04",
   709 => x"f04866c8",
   710 => x"87d0f38e",
   711 => x"5c5b5e0e",
   712 => x"86ec0e5d",
   713 => x"e4c04b71",
   714 => x"28c94866",
   715 => x"c258a6c8",
   716 => x"4abfd6ed",
   717 => x"4872baff",
   718 => x"cc9866c4",
   719 => x"9b7358a6",
   720 => x"87c2c302",
   721 => x"6949a3c8",
   722 => x"87fac202",
   723 => x"986b4872",
   724 => x"c458a6d0",
   725 => x"7e6c4ca3",
   726 => x"cc4866c8",
   727 => x"c605a866",
   728 => x"7b66c487",
   729 => x"c887cdc2",
   730 => x"49731e66",
   731 => x"c487fcfb",
   732 => x"c04d7086",
   733 => x"d004adb7",
   734 => x"4aa3d487",
   735 => x"91c84975",
   736 => x"2149a172",
   737 => x"c77c697b",
   738 => x"cc7bc087",
   739 => x"7c6949a3",
   740 => x"6b4866c4",
   741 => x"58a6c888",
   742 => x"731e66cc",
   743 => x"87cbfb49",
   744 => x"4d7086c4",
   745 => x"49a3c4c1",
   746 => x"6948a6d0",
   747 => x"4866cc78",
   748 => x"06a866d0",
   749 => x"c087f2c0",
   750 => x"c004adb7",
   751 => x"a6c887eb",
   752 => x"78a3d448",
   753 => x"91c84975",
   754 => x"cc8166c8",
   755 => x"88694866",
   756 => x"66d04970",
   757 => x"87d106a9",
   758 => x"dafb4973",
   759 => x"c8497087",
   760 => x"8166c891",
   761 => x"6e4166cc",
   762 => x"4966c479",
   763 => x"f649731e",
   764 => x"86c487c1",
   765 => x"1ed2e5c2",
   766 => x"d0f74973",
   767 => x"d086c487",
   768 => x"e4c049a3",
   769 => x"8eec7966",
   770 => x"1e87e1ef",
   771 => x"4b711e73",
   772 => x"e4c0029b",
   773 => x"fff1c287",
   774 => x"c24a735b",
   775 => x"d2edc28a",
   776 => x"c29249bf",
   777 => x"48bfebf1",
   778 => x"f2c28072",
   779 => x"487158c3",
   780 => x"edc230c4",
   781 => x"edc058e2",
   782 => x"fbf1c287",
   783 => x"eff1c248",
   784 => x"f1c278bf",
   785 => x"f1c248ff",
   786 => x"c278bff3",
   787 => x"02bfdaed",
   788 => x"edc287c9",
   789 => x"c449bfd2",
   790 => x"c287c731",
   791 => x"49bff7f1",
   792 => x"edc231c4",
   793 => x"c7ee59e2",
   794 => x"5b5e0e87",
   795 => x"4a710e5c",
   796 => x"9a724bc0",
   797 => x"87e1c002",
   798 => x"9f49a2da",
   799 => x"edc24b69",
   800 => x"cf02bfda",
   801 => x"49a2d487",
   802 => x"4c49699f",
   803 => x"9cffffc0",
   804 => x"87c234d0",
   805 => x"49744cc0",
   806 => x"fd4973b3",
   807 => x"cded87ed",
   808 => x"5b5e0e87",
   809 => x"f40e5d5c",
   810 => x"c04a7186",
   811 => x"029a727e",
   812 => x"e5c287d8",
   813 => x"78c048ce",
   814 => x"48c6e5c2",
   815 => x"bffff1c2",
   816 => x"cae5c278",
   817 => x"fbf1c248",
   818 => x"edc278bf",
   819 => x"50c048ef",
   820 => x"bfdeedc2",
   821 => x"cee5c249",
   822 => x"aa714abf",
   823 => x"87cac403",
   824 => x"99cf4972",
   825 => x"87eac005",
   826 => x"48fdf9c0",
   827 => x"bfc6e5c2",
   828 => x"d2e5c278",
   829 => x"c6e5c21e",
   830 => x"e5c249bf",
   831 => x"a1c148c6",
   832 => x"ddff7178",
   833 => x"86c487e8",
   834 => x"48f9f9c0",
   835 => x"78d2e5c2",
   836 => x"f9c087cc",
   837 => x"c048bff9",
   838 => x"f9c080e0",
   839 => x"e5c258fd",
   840 => x"c148bfce",
   841 => x"d2e5c280",
   842 => x"0e792758",
   843 => x"97bf0000",
   844 => x"029d4dbf",
   845 => x"c387e3c2",
   846 => x"c202ade5",
   847 => x"f9c087dc",
   848 => x"cb4bbff9",
   849 => x"4c1149a3",
   850 => x"c105accf",
   851 => x"497587d2",
   852 => x"89c199df",
   853 => x"edc291cd",
   854 => x"a3c181e2",
   855 => x"c351124a",
   856 => x"51124aa3",
   857 => x"124aa3c5",
   858 => x"4aa3c751",
   859 => x"a3c95112",
   860 => x"ce51124a",
   861 => x"51124aa3",
   862 => x"124aa3d0",
   863 => x"4aa3d251",
   864 => x"a3d45112",
   865 => x"d651124a",
   866 => x"51124aa3",
   867 => x"124aa3d8",
   868 => x"4aa3dc51",
   869 => x"a3de5112",
   870 => x"c151124a",
   871 => x"87fac07e",
   872 => x"99c84974",
   873 => x"87ebc005",
   874 => x"99d04974",
   875 => x"dc87d105",
   876 => x"cbc00266",
   877 => x"dc497387",
   878 => x"98700f66",
   879 => x"87d3c002",
   880 => x"c6c0056e",
   881 => x"e2edc287",
   882 => x"c050c048",
   883 => x"48bff9f9",
   884 => x"c287e1c2",
   885 => x"c048efed",
   886 => x"edc27e50",
   887 => x"c249bfde",
   888 => x"4abfcee5",
   889 => x"fb04aa71",
   890 => x"f1c287f6",
   891 => x"c005bfff",
   892 => x"edc287c8",
   893 => x"c102bfda",
   894 => x"e5c287f8",
   895 => x"e749bfca",
   896 => x"497087f2",
   897 => x"59cee5c2",
   898 => x"c248a6c4",
   899 => x"78bfcae5",
   900 => x"bfdaedc2",
   901 => x"87d8c002",
   902 => x"cf4966c4",
   903 => x"f8ffffff",
   904 => x"c002a999",
   905 => x"4cc087c5",
   906 => x"c187e1c0",
   907 => x"87dcc04c",
   908 => x"cf4966c4",
   909 => x"a999f8ff",
   910 => x"87c8c002",
   911 => x"c048a6c8",
   912 => x"87c5c078",
   913 => x"c148a6c8",
   914 => x"4c66c878",
   915 => x"c0059c74",
   916 => x"66c487e0",
   917 => x"c289c249",
   918 => x"4abfd2ed",
   919 => x"ebf1c291",
   920 => x"e5c24abf",
   921 => x"a17248c6",
   922 => x"cee5c278",
   923 => x"f978c048",
   924 => x"48c087de",
   925 => x"f3e58ef4",
   926 => x"00000087",
   927 => x"ffffff00",
   928 => x"000e89ff",
   929 => x"000e9200",
   930 => x"54414600",
   931 => x"20203233",
   932 => x"41460020",
   933 => x"20363154",
   934 => x"1e002020",
   935 => x"c348d4ff",
   936 => x"486878ff",
   937 => x"ff1e4f26",
   938 => x"ffc348d4",
   939 => x"48d0ff78",
   940 => x"ff78e1c0",
   941 => x"78d448d4",
   942 => x"48c3f2c2",
   943 => x"50bfd4ff",
   944 => x"ff1e4f26",
   945 => x"e0c048d0",
   946 => x"1e4f2678",
   947 => x"7087ccff",
   948 => x"c6029949",
   949 => x"a9fbc087",
   950 => x"7187f105",
   951 => x"0e4f2648",
   952 => x"0e5c5b5e",
   953 => x"4cc04b71",
   954 => x"7087f0fe",
   955 => x"c0029949",
   956 => x"ecc087f9",
   957 => x"f2c002a9",
   958 => x"a9fbc087",
   959 => x"87ebc002",
   960 => x"acb766cc",
   961 => x"d087c703",
   962 => x"87c20266",
   963 => x"99715371",
   964 => x"c187c202",
   965 => x"87c3fe84",
   966 => x"02994970",
   967 => x"ecc087cd",
   968 => x"87c702a9",
   969 => x"05a9fbc0",
   970 => x"d087d5ff",
   971 => x"87c30266",
   972 => x"c07b97c0",
   973 => x"c405a9ec",
   974 => x"c54a7487",
   975 => x"c04a7487",
   976 => x"48728a0a",
   977 => x"4d2687c2",
   978 => x"4b264c26",
   979 => x"fd1e4f26",
   980 => x"497087c9",
   981 => x"aaf0c04a",
   982 => x"c087c904",
   983 => x"c301aaf9",
   984 => x"8af0c087",
   985 => x"04aac1c1",
   986 => x"dac187c9",
   987 => x"87c301aa",
   988 => x"728af7c0",
   989 => x"0e4f2648",
   990 => x"0e5c5b5e",
   991 => x"d4ff4a71",
   992 => x"c049724c",
   993 => x"4b7087e9",
   994 => x"87c2029b",
   995 => x"d0ff8bc1",
   996 => x"c178c548",
   997 => x"49737cd5",
   998 => x"eac131c6",
   999 => x"4abf97e9",
  1000 => x"70b07148",
  1001 => x"48d0ff7c",
  1002 => x"487378c4",
  1003 => x"0e87d9fe",
  1004 => x"5d5c5b5e",
  1005 => x"7186f80e",
  1006 => x"fb7ec04c",
  1007 => x"4bc087e8",
  1008 => x"97dcc1c1",
  1009 => x"a9c049bf",
  1010 => x"fb87cf04",
  1011 => x"83c187fd",
  1012 => x"97dcc1c1",
  1013 => x"06ab49bf",
  1014 => x"c1c187f1",
  1015 => x"02bf97dc",
  1016 => x"f6fa87cf",
  1017 => x"99497087",
  1018 => x"c087c602",
  1019 => x"f105a9ec",
  1020 => x"fa4bc087",
  1021 => x"4d7087e5",
  1022 => x"c887e0fa",
  1023 => x"dafa58a6",
  1024 => x"c14a7087",
  1025 => x"49a4c883",
  1026 => x"ad496997",
  1027 => x"c087c702",
  1028 => x"c005adff",
  1029 => x"a4c987e7",
  1030 => x"49699749",
  1031 => x"02a966c4",
  1032 => x"c04887c7",
  1033 => x"d405a8ff",
  1034 => x"49a4ca87",
  1035 => x"aa496997",
  1036 => x"c087c602",
  1037 => x"c405aaff",
  1038 => x"d07ec187",
  1039 => x"adecc087",
  1040 => x"c087c602",
  1041 => x"c405adfb",
  1042 => x"c14bc087",
  1043 => x"fe026e7e",
  1044 => x"edf987e1",
  1045 => x"f8487387",
  1046 => x"87eafb8e",
  1047 => x"5b5e0e00",
  1048 => x"f80e5d5c",
  1049 => x"ff4d7186",
  1050 => x"1e754bd4",
  1051 => x"49c8f2c2",
  1052 => x"87f2dfff",
  1053 => x"987086c4",
  1054 => x"87ccc402",
  1055 => x"c148a6c4",
  1056 => x"78bfebea",
  1057 => x"eefb4975",
  1058 => x"48d0ff87",
  1059 => x"d6c178c5",
  1060 => x"754ac07b",
  1061 => x"7b1149a2",
  1062 => x"b7cb82c1",
  1063 => x"87f304aa",
  1064 => x"ffc34acc",
  1065 => x"c082c17b",
  1066 => x"04aab7e0",
  1067 => x"d0ff87f4",
  1068 => x"c378c448",
  1069 => x"78c57bff",
  1070 => x"c17bd3c1",
  1071 => x"6678c47b",
  1072 => x"a8b7c048",
  1073 => x"87f0c206",
  1074 => x"bfd0f2c2",
  1075 => x"4866c44c",
  1076 => x"a6c88874",
  1077 => x"029c7458",
  1078 => x"c287f9c1",
  1079 => x"c87ed2e5",
  1080 => x"c08c4dc0",
  1081 => x"c603acb7",
  1082 => x"a4c0c887",
  1083 => x"c24cc04d",
  1084 => x"bf97c3f2",
  1085 => x"0299d049",
  1086 => x"1ec087d1",
  1087 => x"49c8f2c2",
  1088 => x"c487cae3",
  1089 => x"4a497086",
  1090 => x"c287eec0",
  1091 => x"c21ed2e5",
  1092 => x"e249c8f2",
  1093 => x"86c487f7",
  1094 => x"ff4a4970",
  1095 => x"c5c848d0",
  1096 => x"7bd4c178",
  1097 => x"7bbf976e",
  1098 => x"80c1486e",
  1099 => x"8dc17e70",
  1100 => x"87f0ff05",
  1101 => x"c448d0ff",
  1102 => x"059a7278",
  1103 => x"48c087c5",
  1104 => x"c187c7c1",
  1105 => x"c8f2c21e",
  1106 => x"87e7e049",
  1107 => x"9c7486c4",
  1108 => x"87c7fe05",
  1109 => x"c04866c4",
  1110 => x"d106a8b7",
  1111 => x"c8f2c287",
  1112 => x"d078c048",
  1113 => x"f478c080",
  1114 => x"d4f2c280",
  1115 => x"66c478bf",
  1116 => x"a8b7c048",
  1117 => x"87d0fd01",
  1118 => x"c548d0ff",
  1119 => x"7bd3c178",
  1120 => x"78c47bc0",
  1121 => x"87c248c1",
  1122 => x"8ef848c0",
  1123 => x"4c264d26",
  1124 => x"4f264b26",
  1125 => x"5c5b5e0e",
  1126 => x"711e0e5d",
  1127 => x"4d4cc04b",
  1128 => x"e8c004ab",
  1129 => x"effec087",
  1130 => x"029d751e",
  1131 => x"4ac087c4",
  1132 => x"4ac187c2",
  1133 => x"e8eb4972",
  1134 => x"7086c487",
  1135 => x"6e84c17e",
  1136 => x"7387c205",
  1137 => x"7385c14c",
  1138 => x"d8ff06ac",
  1139 => x"26486e87",
  1140 => x"0e87f9fe",
  1141 => x"0e5c5b5e",
  1142 => x"66cc4b71",
  1143 => x"4c87d802",
  1144 => x"028cf0c0",
  1145 => x"4a7487d8",
  1146 => x"d1028ac1",
  1147 => x"cd028a87",
  1148 => x"c9028a87",
  1149 => x"7387d987",
  1150 => x"87e1f949",
  1151 => x"1e7487d2",
  1152 => x"d8c149c0",
  1153 => x"1e7487fb",
  1154 => x"d8c14973",
  1155 => x"86c887f3",
  1156 => x"0e87fbfd",
  1157 => x"5d5c5b5e",
  1158 => x"4c711e0e",
  1159 => x"c291de49",
  1160 => x"714de4f3",
  1161 => x"026d9785",
  1162 => x"c287dcc1",
  1163 => x"4abfd0f3",
  1164 => x"49728274",
  1165 => x"7087ddfd",
  1166 => x"c0026e7e",
  1167 => x"f3c287f2",
  1168 => x"4a6e4bd8",
  1169 => x"f9fe49cb",
  1170 => x"4b7487de",
  1171 => x"eac193cb",
  1172 => x"83c483fd",
  1173 => x"7bcbcac1",
  1174 => x"c1c14974",
  1175 => x"7b7587f0",
  1176 => x"97eaeac1",
  1177 => x"c21e49bf",
  1178 => x"fd49d8f3",
  1179 => x"86c487e5",
  1180 => x"c1c14974",
  1181 => x"49c087d8",
  1182 => x"87f7c2c1",
  1183 => x"48c4f2c2",
  1184 => x"49c178c0",
  1185 => x"2687dadd",
  1186 => x"4c87c1fc",
  1187 => x"6964616f",
  1188 => x"2e2e676e",
  1189 => x"5e0e002e",
  1190 => x"710e5c5b",
  1191 => x"f3c24a4b",
  1192 => x"7282bfd0",
  1193 => x"87ecfb49",
  1194 => x"029c4c70",
  1195 => x"e64987c4",
  1196 => x"f3c287f7",
  1197 => x"78c048d0",
  1198 => x"e4dc49c1",
  1199 => x"87cefb87",
  1200 => x"5c5b5e0e",
  1201 => x"86f40e5d",
  1202 => x"4dd2e5c2",
  1203 => x"a6c44cc0",
  1204 => x"c278c048",
  1205 => x"49bfd0f3",
  1206 => x"c106a9c0",
  1207 => x"e5c287c1",
  1208 => x"029848d2",
  1209 => x"c087f8c0",
  1210 => x"c81eeffe",
  1211 => x"87c70266",
  1212 => x"c048a6c4",
  1213 => x"c487c578",
  1214 => x"78c148a6",
  1215 => x"e64966c4",
  1216 => x"86c487df",
  1217 => x"84c14d70",
  1218 => x"c14866c4",
  1219 => x"58a6c880",
  1220 => x"bfd0f3c2",
  1221 => x"c603ac49",
  1222 => x"059d7587",
  1223 => x"c087c8ff",
  1224 => x"029d754c",
  1225 => x"c087e0c3",
  1226 => x"c81eeffe",
  1227 => x"87c70266",
  1228 => x"c048a6cc",
  1229 => x"cc87c578",
  1230 => x"78c148a6",
  1231 => x"e54966cc",
  1232 => x"86c487df",
  1233 => x"026e7e70",
  1234 => x"6e87e9c2",
  1235 => x"9781cb49",
  1236 => x"99d04969",
  1237 => x"87d6c102",
  1238 => x"4ad6cac1",
  1239 => x"91cb4974",
  1240 => x"81fdeac1",
  1241 => x"81c87972",
  1242 => x"7451ffc3",
  1243 => x"c291de49",
  1244 => x"714de4f3",
  1245 => x"97c1c285",
  1246 => x"49a5c17d",
  1247 => x"c251e0c0",
  1248 => x"bf97e2ed",
  1249 => x"c187d202",
  1250 => x"4ba5c284",
  1251 => x"4ae2edc2",
  1252 => x"f4fe49db",
  1253 => x"dbc187d2",
  1254 => x"49a5cd87",
  1255 => x"84c151c0",
  1256 => x"6e4ba5c2",
  1257 => x"fe49cb4a",
  1258 => x"c187fdf3",
  1259 => x"c8c187c6",
  1260 => x"49744ad3",
  1261 => x"eac191cb",
  1262 => x"797281fd",
  1263 => x"97e2edc2",
  1264 => x"87d802bf",
  1265 => x"91de4974",
  1266 => x"f3c284c1",
  1267 => x"83714be4",
  1268 => x"4ae2edc2",
  1269 => x"f3fe49dd",
  1270 => x"87d887ce",
  1271 => x"93de4b74",
  1272 => x"83e4f3c2",
  1273 => x"c049a3cb",
  1274 => x"7384c151",
  1275 => x"49cb4a6e",
  1276 => x"87f4f2fe",
  1277 => x"c14866c4",
  1278 => x"58a6c880",
  1279 => x"c003acc7",
  1280 => x"056e87c5",
  1281 => x"7487e0fc",
  1282 => x"f58ef448",
  1283 => x"731e87fe",
  1284 => x"494b711e",
  1285 => x"eac191cb",
  1286 => x"a1c881fd",
  1287 => x"e9eac14a",
  1288 => x"c9501248",
  1289 => x"c1c14aa1",
  1290 => x"501248dc",
  1291 => x"eac181ca",
  1292 => x"501148ea",
  1293 => x"97eaeac1",
  1294 => x"c01e49bf",
  1295 => x"87d3f649",
  1296 => x"48c4f2c2",
  1297 => x"49c178de",
  1298 => x"2687d6d6",
  1299 => x"1e87c1f5",
  1300 => x"cb494a71",
  1301 => x"fdeac191",
  1302 => x"1181c881",
  1303 => x"c8f2c248",
  1304 => x"d0f3c258",
  1305 => x"c178c048",
  1306 => x"87f5d549",
  1307 => x"c01e4f26",
  1308 => x"fefac049",
  1309 => x"1e4f2687",
  1310 => x"d2029971",
  1311 => x"d2ecc187",
  1312 => x"f750c048",
  1313 => x"cfd1c180",
  1314 => x"f6eac140",
  1315 => x"c187ce78",
  1316 => x"c148ceec",
  1317 => x"fc78efea",
  1318 => x"eed1c180",
  1319 => x"0e4f2678",
  1320 => x"0e5c5b5e",
  1321 => x"cb4a4c71",
  1322 => x"fdeac192",
  1323 => x"49a2c882",
  1324 => x"974ba2c9",
  1325 => x"971e4b6b",
  1326 => x"ca1e4969",
  1327 => x"c0491282",
  1328 => x"c087f9e5",
  1329 => x"87d9d449",
  1330 => x"f8c04974",
  1331 => x"8ef887c0",
  1332 => x"1e87fbf2",
  1333 => x"4b711e73",
  1334 => x"87c3ff49",
  1335 => x"fefe4973",
  1336 => x"87ecf287",
  1337 => x"711e731e",
  1338 => x"4aa3c64b",
  1339 => x"c187db02",
  1340 => x"87d6028a",
  1341 => x"dac1028a",
  1342 => x"c0028a87",
  1343 => x"028a87fc",
  1344 => x"8a87e1c0",
  1345 => x"c187cb02",
  1346 => x"49c787db",
  1347 => x"c187c0fd",
  1348 => x"f3c287de",
  1349 => x"c102bfd0",
  1350 => x"c14887cb",
  1351 => x"d4f3c288",
  1352 => x"87c1c158",
  1353 => x"bfd4f3c2",
  1354 => x"87f9c002",
  1355 => x"bfd0f3c2",
  1356 => x"c280c148",
  1357 => x"c058d4f3",
  1358 => x"f3c287eb",
  1359 => x"c649bfd0",
  1360 => x"d4f3c289",
  1361 => x"a9b7c059",
  1362 => x"c287da03",
  1363 => x"c048d0f3",
  1364 => x"c287d278",
  1365 => x"02bfd4f3",
  1366 => x"f3c287cb",
  1367 => x"c648bfd0",
  1368 => x"d4f3c280",
  1369 => x"d149c058",
  1370 => x"497387f7",
  1371 => x"87def5c0",
  1372 => x"0e87ddf0",
  1373 => x"5d5c5b5e",
  1374 => x"86d0ff0e",
  1375 => x"c859a6dc",
  1376 => x"78c048a6",
  1377 => x"c4c180c4",
  1378 => x"80c47866",
  1379 => x"80c478c1",
  1380 => x"f3c278c1",
  1381 => x"78c148d4",
  1382 => x"bfc4f2c2",
  1383 => x"05a8de48",
  1384 => x"dbf487cb",
  1385 => x"cc497087",
  1386 => x"f3cf59a6",
  1387 => x"87f6e387",
  1388 => x"e387d8e4",
  1389 => x"4c7087e5",
  1390 => x"02acfbc0",
  1391 => x"d887fbc1",
  1392 => x"edc10566",
  1393 => x"66c0c187",
  1394 => x"6a82c44a",
  1395 => x"c11e727e",
  1396 => x"c448d5e7",
  1397 => x"a1c84966",
  1398 => x"7141204a",
  1399 => x"87f905aa",
  1400 => x"4a265110",
  1401 => x"4866c0c1",
  1402 => x"78ced0c1",
  1403 => x"81c7496a",
  1404 => x"c0c15174",
  1405 => x"81c84966",
  1406 => x"c0c151c1",
  1407 => x"81c94966",
  1408 => x"c0c151c0",
  1409 => x"81ca4966",
  1410 => x"1ec151c0",
  1411 => x"496a1ed8",
  1412 => x"cae381c8",
  1413 => x"c186c887",
  1414 => x"c04866c4",
  1415 => x"87c701a8",
  1416 => x"c148a6c8",
  1417 => x"c187ce78",
  1418 => x"c14866c4",
  1419 => x"58a6d088",
  1420 => x"d6e287c3",
  1421 => x"48a6d087",
  1422 => x"9c7478c2",
  1423 => x"87dccd02",
  1424 => x"c14866c8",
  1425 => x"03a866c8",
  1426 => x"dc87d1cd",
  1427 => x"78c048a6",
  1428 => x"78c080e8",
  1429 => x"7087c4e1",
  1430 => x"acd0c14c",
  1431 => x"87d8c205",
  1432 => x"e37e66c4",
  1433 => x"497087e8",
  1434 => x"e059a6c8",
  1435 => x"4c7087ed",
  1436 => x"05acecc0",
  1437 => x"c887ecc1",
  1438 => x"91cb4966",
  1439 => x"8166c0c1",
  1440 => x"6a4aa1c4",
  1441 => x"4aa1c84d",
  1442 => x"c15266c4",
  1443 => x"e079cfd1",
  1444 => x"4c7087c9",
  1445 => x"87d9029c",
  1446 => x"02acfbc0",
  1447 => x"557487d3",
  1448 => x"87f7dfff",
  1449 => x"029c4c70",
  1450 => x"fbc087c7",
  1451 => x"edff05ac",
  1452 => x"55e0c087",
  1453 => x"c055c1c2",
  1454 => x"66d87d97",
  1455 => x"05a96e49",
  1456 => x"66c887db",
  1457 => x"a866cc48",
  1458 => x"c887ca04",
  1459 => x"80c14866",
  1460 => x"c858a6cc",
  1461 => x"4866cc87",
  1462 => x"a6d088c1",
  1463 => x"fadeff58",
  1464 => x"c14c7087",
  1465 => x"c805acd0",
  1466 => x"4866d487",
  1467 => x"a6d880c1",
  1468 => x"acd0c158",
  1469 => x"87e8fd02",
  1470 => x"48a6e0c0",
  1471 => x"c47866d8",
  1472 => x"e0c04866",
  1473 => x"c905a866",
  1474 => x"e4c087e4",
  1475 => x"78c048a6",
  1476 => x"78c080c4",
  1477 => x"fbc04874",
  1478 => x"6e7e7088",
  1479 => x"87e7c802",
  1480 => x"88cb486e",
  1481 => x"026e7e70",
  1482 => x"6e87cdc1",
  1483 => x"7088c948",
  1484 => x"c3026e7e",
  1485 => x"486e87e9",
  1486 => x"7e7088c4",
  1487 => x"87ce026e",
  1488 => x"88c1486e",
  1489 => x"026e7e70",
  1490 => x"c787d4c3",
  1491 => x"a6dc87f3",
  1492 => x"78f0c048",
  1493 => x"87c3ddff",
  1494 => x"ecc04c70",
  1495 => x"c4c002ac",
  1496 => x"a6e0c087",
  1497 => x"acecc05c",
  1498 => x"ff87cd02",
  1499 => x"7087ecdc",
  1500 => x"acecc04c",
  1501 => x"87f3ff05",
  1502 => x"02acecc0",
  1503 => x"ff87c4c0",
  1504 => x"c087d8dc",
  1505 => x"d01eca1e",
  1506 => x"91cb4966",
  1507 => x"4866c8c1",
  1508 => x"a6cc8071",
  1509 => x"4866c858",
  1510 => x"a6d080c4",
  1511 => x"bf66cc58",
  1512 => x"fadcff49",
  1513 => x"de1ec187",
  1514 => x"bf66d41e",
  1515 => x"eedcff49",
  1516 => x"7086d087",
  1517 => x"8909c049",
  1518 => x"59a6ecc0",
  1519 => x"4866e8c0",
  1520 => x"c006a8c0",
  1521 => x"e8c087ee",
  1522 => x"a8dd4866",
  1523 => x"87e4c003",
  1524 => x"49bf66c4",
  1525 => x"8166e8c0",
  1526 => x"c051e0c0",
  1527 => x"c14966e8",
  1528 => x"bf66c481",
  1529 => x"51c1c281",
  1530 => x"4966e8c0",
  1531 => x"66c481c2",
  1532 => x"51c081bf",
  1533 => x"d0c1486e",
  1534 => x"496e78ce",
  1535 => x"66d081c8",
  1536 => x"c9496e51",
  1537 => x"5166d481",
  1538 => x"81ca496e",
  1539 => x"d05166dc",
  1540 => x"80c14866",
  1541 => x"4858a6d4",
  1542 => x"78c180d8",
  1543 => x"ff87e8c4",
  1544 => x"7087ebdc",
  1545 => x"a6ecc049",
  1546 => x"e1dcff59",
  1547 => x"c0497087",
  1548 => x"dc59a6e0",
  1549 => x"ecc04866",
  1550 => x"cac005a8",
  1551 => x"48a6dc87",
  1552 => x"7866e8c0",
  1553 => x"ff87c4c0",
  1554 => x"c887d0d9",
  1555 => x"91cb4966",
  1556 => x"4866c0c1",
  1557 => x"7e708071",
  1558 => x"82c84a6e",
  1559 => x"81ca496e",
  1560 => x"5166e8c0",
  1561 => x"c14966dc",
  1562 => x"66e8c081",
  1563 => x"7148c189",
  1564 => x"c1497030",
  1565 => x"7a977189",
  1566 => x"bfc0f7c2",
  1567 => x"66e8c049",
  1568 => x"4a6a9729",
  1569 => x"c0987148",
  1570 => x"6e58a6f0",
  1571 => x"6981c449",
  1572 => x"66e0c04d",
  1573 => x"a866c448",
  1574 => x"87c8c002",
  1575 => x"c048a6c4",
  1576 => x"87c5c078",
  1577 => x"c148a6c4",
  1578 => x"1e66c478",
  1579 => x"751ee0c0",
  1580 => x"ead8ff49",
  1581 => x"7086c887",
  1582 => x"acb7c04c",
  1583 => x"87d4c106",
  1584 => x"e0c08574",
  1585 => x"75897449",
  1586 => x"dee7c14b",
  1587 => x"dffe714a",
  1588 => x"85c287d6",
  1589 => x"4866e4c0",
  1590 => x"e8c080c1",
  1591 => x"ecc058a6",
  1592 => x"81c14966",
  1593 => x"c002a970",
  1594 => x"a6c487c8",
  1595 => x"c078c048",
  1596 => x"a6c487c5",
  1597 => x"c478c148",
  1598 => x"a4c21e66",
  1599 => x"48e0c049",
  1600 => x"49708871",
  1601 => x"ff49751e",
  1602 => x"c887d4d7",
  1603 => x"a8b7c086",
  1604 => x"87c0ff01",
  1605 => x"0266e4c0",
  1606 => x"6e87d1c0",
  1607 => x"c081c949",
  1608 => x"6e5166e4",
  1609 => x"dfd2c148",
  1610 => x"87ccc078",
  1611 => x"81c9496e",
  1612 => x"486e51c2",
  1613 => x"78d3d3c1",
  1614 => x"48a6e8c0",
  1615 => x"c6c078c1",
  1616 => x"c6d6ff87",
  1617 => x"c04c7087",
  1618 => x"c00266e8",
  1619 => x"66c887f5",
  1620 => x"a866cc48",
  1621 => x"87cbc004",
  1622 => x"c14866c8",
  1623 => x"58a6cc80",
  1624 => x"cc87e0c0",
  1625 => x"88c14866",
  1626 => x"c058a6d0",
  1627 => x"c6c187d5",
  1628 => x"c8c005ac",
  1629 => x"4866d087",
  1630 => x"a6d480c1",
  1631 => x"cad5ff58",
  1632 => x"d44c7087",
  1633 => x"80c14866",
  1634 => x"7458a6d8",
  1635 => x"cbc0029c",
  1636 => x"4866c887",
  1637 => x"a866c8c1",
  1638 => x"87eff204",
  1639 => x"87e2d4ff",
  1640 => x"c74866c8",
  1641 => x"e5c003a8",
  1642 => x"d4f3c287",
  1643 => x"c878c048",
  1644 => x"91cb4966",
  1645 => x"8166c0c1",
  1646 => x"6a4aa1c4",
  1647 => x"7952c04a",
  1648 => x"c14866c8",
  1649 => x"58a6cc80",
  1650 => x"ff04a8c7",
  1651 => x"d0ff87db",
  1652 => x"f7deff8e",
  1653 => x"616f4c87",
  1654 => x"2e2a2064",
  1655 => x"203a0020",
  1656 => x"1e731e00",
  1657 => x"029b4b71",
  1658 => x"f3c287c6",
  1659 => x"78c048d0",
  1660 => x"f3c21ec7",
  1661 => x"1e49bfd0",
  1662 => x"1efdeac1",
  1663 => x"bfc4f2c2",
  1664 => x"87efed49",
  1665 => x"f2c286cc",
  1666 => x"e949bfc4",
  1667 => x"9b7387e9",
  1668 => x"c187c802",
  1669 => x"c049fdea",
  1670 => x"ff87c5e4",
  1671 => x"1e87f1dd",
  1672 => x"c187d4c7",
  1673 => x"87f9fe49",
  1674 => x"87c9e4fe",
  1675 => x"cd029870",
  1676 => x"c4edfe87",
  1677 => x"02987087",
  1678 => x"4ac187c4",
  1679 => x"4ac087c2",
  1680 => x"ce059a72",
  1681 => x"c11ec087",
  1682 => x"c049f0e9",
  1683 => x"c487d7f0",
  1684 => x"c087fe86",
  1685 => x"fbe9c11e",
  1686 => x"c9f0c049",
  1687 => x"c01ec087",
  1688 => x"7087cdfa",
  1689 => x"fdefc049",
  1690 => x"87cac387",
  1691 => x"4f268ef8",
  1692 => x"66204453",
  1693 => x"656c6961",
  1694 => x"42002e64",
  1695 => x"69746f6f",
  1696 => x"2e2e676e",
  1697 => x"c01e002e",
  1698 => x"c087f1e6",
  1699 => x"f687def3",
  1700 => x"1e4f2687",
  1701 => x"48d0f3c2",
  1702 => x"f2c278c0",
  1703 => x"78c048c4",
  1704 => x"e187fcfd",
  1705 => x"2648c087",
  1706 => x"0100004f",
  1707 => x"80000000",
  1708 => x"69784520",
  1709 => x"20800074",
  1710 => x"6b636142",
  1711 => x"00121300",
  1712 => x"002ce400",
  1713 => x"00000000",
  1714 => x"00001213",
  1715 => x"00002d02",
  1716 => x"13000000",
  1717 => x"20000012",
  1718 => x"0000002d",
  1719 => x"12130000",
  1720 => x"2d3e0000",
  1721 => x"00000000",
  1722 => x"00121300",
  1723 => x"002d5c00",
  1724 => x"00000000",
  1725 => x"00001213",
  1726 => x"00002d7a",
  1727 => x"13000000",
  1728 => x"98000012",
  1729 => x"0000002d",
  1730 => x"144f0000",
  1731 => x"00000000",
  1732 => x"00000000",
  1733 => x"0014e400",
  1734 => x"00000000",
  1735 => x"00000000",
  1736 => x"48f0fe1e",
  1737 => x"09cd78c0",
  1738 => x"4f260979",
  1739 => x"f0fe1e1e",
  1740 => x"26487ebf",
  1741 => x"fe1e4f26",
  1742 => x"78c148f0",
  1743 => x"fe1e4f26",
  1744 => x"78c048f0",
  1745 => x"711e4f26",
  1746 => x"5252c04a",
  1747 => x"5e0e4f26",
  1748 => x"0e5d5c5b",
  1749 => x"4d7186f4",
  1750 => x"c17e6d97",
  1751 => x"6c974ca5",
  1752 => x"58a6c848",
  1753 => x"66c4486e",
  1754 => x"87c505a8",
  1755 => x"e6c048ff",
  1756 => x"87caff87",
  1757 => x"9749a5c2",
  1758 => x"a3714b6c",
  1759 => x"4b6b974b",
  1760 => x"6e7e6c97",
  1761 => x"c880c148",
  1762 => x"98c758a6",
  1763 => x"7058a6cc",
  1764 => x"e1fe7c97",
  1765 => x"f4487387",
  1766 => x"264d268e",
  1767 => x"264b264c",
  1768 => x"5b5e0e4f",
  1769 => x"86f40e5c",
  1770 => x"66d84c71",
  1771 => x"9affc34a",
  1772 => x"974ba4c2",
  1773 => x"a173496c",
  1774 => x"97517249",
  1775 => x"486e7e6c",
  1776 => x"a6c880c1",
  1777 => x"cc98c758",
  1778 => x"547058a6",
  1779 => x"caff8ef4",
  1780 => x"fd1e1e87",
  1781 => x"bfe087e8",
  1782 => x"e0c0494a",
  1783 => x"cb0299c0",
  1784 => x"c21e7287",
  1785 => x"fe49f6f6",
  1786 => x"86c487f7",
  1787 => x"7087fdfc",
  1788 => x"87c2fd7e",
  1789 => x"1e4f2626",
  1790 => x"49f6f6c2",
  1791 => x"c187c7fd",
  1792 => x"fc49d1ef",
  1793 => x"f7c387da",
  1794 => x"0e4f2687",
  1795 => x"5d5c5b5e",
  1796 => x"c24d710e",
  1797 => x"fc49f6f6",
  1798 => x"4b7087f4",
  1799 => x"04abb7c0",
  1800 => x"c387c2c3",
  1801 => x"c905abf0",
  1802 => x"eff3c187",
  1803 => x"c278c148",
  1804 => x"e0c387e3",
  1805 => x"87c905ab",
  1806 => x"48f3f3c1",
  1807 => x"d4c278c1",
  1808 => x"f3f3c187",
  1809 => x"87c602bf",
  1810 => x"4ca3c0c2",
  1811 => x"4c7387c2",
  1812 => x"bfeff3c1",
  1813 => x"87e0c002",
  1814 => x"b7c44974",
  1815 => x"f5c19129",
  1816 => x"4a7481cf",
  1817 => x"92c29acf",
  1818 => x"307248c1",
  1819 => x"baff4a70",
  1820 => x"98694872",
  1821 => x"87db7970",
  1822 => x"b7c44974",
  1823 => x"f5c19129",
  1824 => x"4a7481cf",
  1825 => x"92c29acf",
  1826 => x"307248c3",
  1827 => x"69484a70",
  1828 => x"757970b0",
  1829 => x"f0c0059d",
  1830 => x"48d0ff87",
  1831 => x"ff78e1c8",
  1832 => x"78c548d4",
  1833 => x"bff3f3c1",
  1834 => x"c387c302",
  1835 => x"f3c178e0",
  1836 => x"c602bfef",
  1837 => x"48d4ff87",
  1838 => x"ff78f0c3",
  1839 => x"787348d4",
  1840 => x"c848d0ff",
  1841 => x"e0c078e1",
  1842 => x"f3f3c178",
  1843 => x"c178c048",
  1844 => x"c048eff3",
  1845 => x"f6f6c278",
  1846 => x"87f2f949",
  1847 => x"b7c04b70",
  1848 => x"fefc03ab",
  1849 => x"2648c087",
  1850 => x"264c264d",
  1851 => x"004f264b",
  1852 => x"00000000",
  1853 => x"1e000000",
  1854 => x"fc494a71",
  1855 => x"4f2687cd",
  1856 => x"724ac01e",
  1857 => x"c191c449",
  1858 => x"c081cff5",
  1859 => x"d082c179",
  1860 => x"ee04aab7",
  1861 => x"0e4f2687",
  1862 => x"5d5c5b5e",
  1863 => x"f84d710e",
  1864 => x"4a7587dc",
  1865 => x"922ab7c4",
  1866 => x"82cff5c1",
  1867 => x"9ccf4c75",
  1868 => x"496a94c2",
  1869 => x"c32b744b",
  1870 => x"7448c29b",
  1871 => x"ff4c7030",
  1872 => x"714874bc",
  1873 => x"f77a7098",
  1874 => x"487387ec",
  1875 => x"0087d8fe",
  1876 => x"00000000",
  1877 => x"00000000",
  1878 => x"00000000",
  1879 => x"00000000",
  1880 => x"00000000",
  1881 => x"00000000",
  1882 => x"00000000",
  1883 => x"00000000",
  1884 => x"00000000",
  1885 => x"00000000",
  1886 => x"00000000",
  1887 => x"00000000",
  1888 => x"00000000",
  1889 => x"00000000",
  1890 => x"00000000",
  1891 => x"1e000000",
  1892 => x"c848d0ff",
  1893 => x"487178e1",
  1894 => x"7808d4ff",
  1895 => x"ff1e4f26",
  1896 => x"e1c848d0",
  1897 => x"ff487178",
  1898 => x"c47808d4",
  1899 => x"d4ff4866",
  1900 => x"4f267808",
  1901 => x"c44a711e",
  1902 => x"721e4966",
  1903 => x"87deff49",
  1904 => x"c048d0ff",
  1905 => x"262678e0",
  1906 => x"1e731e4f",
  1907 => x"66c84b71",
  1908 => x"4a731e49",
  1909 => x"49a2e0c1",
  1910 => x"2687d9ff",
  1911 => x"4d2687c4",
  1912 => x"4b264c26",
  1913 => x"731e4f26",
  1914 => x"4b4a711e",
  1915 => x"03abb7c2",
  1916 => x"49a387c8",
  1917 => x"9affc34a",
  1918 => x"a3ce87c7",
  1919 => x"ffc34a49",
  1920 => x"4966c89a",
  1921 => x"fe49721e",
  1922 => x"ff2687ea",
  1923 => x"ff1e87d4",
  1924 => x"ffc34ad4",
  1925 => x"48d0ff7a",
  1926 => x"de78e1c0",
  1927 => x"c0f7c27a",
  1928 => x"48497abf",
  1929 => x"7a7028c8",
  1930 => x"28d04871",
  1931 => x"48717a70",
  1932 => x"7a7028d8",
  1933 => x"c048d0ff",
  1934 => x"4f2678e0",
  1935 => x"5c5b5e0e",
  1936 => x"4c710e5d",
  1937 => x"bfc0f7c2",
  1938 => x"2974494d",
  1939 => x"66d04b71",
  1940 => x"d483c19b",
  1941 => x"04abb766",
  1942 => x"4bc087c2",
  1943 => x"744966d0",
  1944 => x"75b9ff31",
  1945 => x"744a7399",
  1946 => x"71487232",
  1947 => x"c4f7c2b0",
  1948 => x"87dafe58",
  1949 => x"4c264d26",
  1950 => x"4f264b26",
  1951 => x"48d0ff1e",
  1952 => x"7178c9c8",
  1953 => x"08d4ff48",
  1954 => x"1e4f2678",
  1955 => x"eb494a71",
  1956 => x"48d0ff87",
  1957 => x"4f2678c8",
  1958 => x"711e731e",
  1959 => x"d0f7c24b",
  1960 => x"87c302bf",
  1961 => x"ff87ebc2",
  1962 => x"c9c848d0",
  1963 => x"c0497378",
  1964 => x"d4ffb1e0",
  1965 => x"c2787148",
  1966 => x"c048c4f7",
  1967 => x"0266c878",
  1968 => x"ffc387c5",
  1969 => x"c087c249",
  1970 => x"ccf7c249",
  1971 => x"0266cc59",
  1972 => x"d5c587c6",
  1973 => x"87c44ad5",
  1974 => x"4affffcf",
  1975 => x"5ad0f7c2",
  1976 => x"48d0f7c2",
  1977 => x"87c478c1",
  1978 => x"4c264d26",
  1979 => x"4f264b26",
  1980 => x"5c5b5e0e",
  1981 => x"4a710e5d",
  1982 => x"bfccf7c2",
  1983 => x"029a724c",
  1984 => x"c84987cb",
  1985 => x"cefac191",
  1986 => x"c483714b",
  1987 => x"cefec187",
  1988 => x"134dc04b",
  1989 => x"c2997449",
  1990 => x"b9bfc8f7",
  1991 => x"7148d4ff",
  1992 => x"2cb7c178",
  1993 => x"adb7c885",
  1994 => x"c287e804",
  1995 => x"48bfc4f7",
  1996 => x"f7c280c8",
  1997 => x"effe58c8",
  1998 => x"1e731e87",
  1999 => x"4a134b71",
  2000 => x"87cb029a",
  2001 => x"e7fe4972",
  2002 => x"9a4a1387",
  2003 => x"fe87f505",
  2004 => x"c21e87da",
  2005 => x"49bfc4f7",
  2006 => x"48c4f7c2",
  2007 => x"c478a1c1",
  2008 => x"03a9b7c0",
  2009 => x"d4ff87db",
  2010 => x"c8f7c248",
  2011 => x"f7c278bf",
  2012 => x"c249bfc4",
  2013 => x"c148c4f7",
  2014 => x"c0c478a1",
  2015 => x"e504a9b7",
  2016 => x"48d0ff87",
  2017 => x"f7c278c8",
  2018 => x"78c048d0",
  2019 => x"00004f26",
  2020 => x"00000000",
  2021 => x"00000000",
  2022 => x"005f5f00",
  2023 => x"03000000",
  2024 => x"03030003",
  2025 => x"7f140000",
  2026 => x"7f7f147f",
  2027 => x"24000014",
  2028 => x"3a6b6b2e",
  2029 => x"6a4c0012",
  2030 => x"566c1836",
  2031 => x"7e300032",
  2032 => x"3a77594f",
  2033 => x"00004068",
  2034 => x"00030704",
  2035 => x"00000000",
  2036 => x"41633e1c",
  2037 => x"00000000",
  2038 => x"1c3e6341",
  2039 => x"2a080000",
  2040 => x"3e1c1c3e",
  2041 => x"0800082a",
  2042 => x"083e3e08",
  2043 => x"00000008",
  2044 => x"0060e080",
  2045 => x"08000000",
  2046 => x"08080808",
  2047 => x"00000008",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
