
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"cc",x"fc",x"c2",x"87"),
    12 => (x"86",x"c0",x"c8",x"4e"),
    13 => (x"49",x"cc",x"fc",x"c2"),
    14 => (x"48",x"ec",x"e4",x"c2"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"c8",x"e9"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"1e",x"73",x"1e",x"72"),
    21 => (x"02",x"11",x"48",x"12"),
    22 => (x"c3",x"4b",x"87",x"ca"),
    23 => (x"73",x"9b",x"98",x"df"),
    24 => (x"87",x"f0",x"02",x"88"),
    25 => (x"4a",x"26",x"4b",x"26"),
    26 => (x"73",x"1e",x"4f",x"26"),
    27 => (x"c1",x"1e",x"72",x"1e"),
    28 => (x"87",x"ca",x"04",x"8b"),
    29 => (x"02",x"11",x"48",x"12"),
    30 => (x"02",x"88",x"87",x"c4"),
    31 => (x"4a",x"26",x"87",x"f1"),
    32 => (x"4f",x"26",x"4b",x"26"),
    33 => (x"73",x"1e",x"74",x"1e"),
    34 => (x"c1",x"1e",x"72",x"1e"),
    35 => (x"87",x"d0",x"04",x"8b"),
    36 => (x"02",x"11",x"48",x"12"),
    37 => (x"c3",x"4c",x"87",x"ca"),
    38 => (x"74",x"9c",x"98",x"df"),
    39 => (x"87",x"eb",x"02",x"88"),
    40 => (x"4b",x"26",x"4a",x"26"),
    41 => (x"4f",x"26",x"4c",x"26"),
    42 => (x"81",x"48",x"73",x"1e"),
    43 => (x"c5",x"02",x"a9",x"73"),
    44 => (x"05",x"53",x"12",x"87"),
    45 => (x"4f",x"26",x"87",x"f6"),
    46 => (x"72",x"1e",x"73",x"1e"),
    47 => (x"e7",x"c0",x"02",x"9a"),
    48 => (x"c1",x"48",x"c0",x"87"),
    49 => (x"06",x"a9",x"72",x"4b"),
    50 => (x"82",x"72",x"87",x"d1"),
    51 => (x"73",x"87",x"c9",x"06"),
    52 => (x"01",x"a9",x"72",x"83"),
    53 => (x"87",x"c3",x"87",x"f4"),
    54 => (x"72",x"3a",x"b2",x"c1"),
    55 => (x"73",x"89",x"03",x"a9"),
    56 => (x"2a",x"c1",x"07",x"80"),
    57 => (x"87",x"f3",x"05",x"2b"),
    58 => (x"4f",x"26",x"4b",x"26"),
    59 => (x"c4",x"1e",x"75",x"1e"),
    60 => (x"a1",x"b7",x"71",x"4d"),
    61 => (x"c1",x"b9",x"ff",x"04"),
    62 => (x"07",x"bd",x"c3",x"81"),
    63 => (x"04",x"a2",x"b7",x"72"),
    64 => (x"82",x"c1",x"ba",x"ff"),
    65 => (x"fe",x"07",x"bd",x"c1"),
    66 => (x"2d",x"c1",x"87",x"ee"),
    67 => (x"c1",x"b8",x"ff",x"04"),
    68 => (x"04",x"2d",x"07",x"80"),
    69 => (x"81",x"c1",x"b9",x"ff"),
    70 => (x"26",x"4d",x"26",x"07"),
    71 => (x"4a",x"71",x"1e",x"4f"),
    72 => (x"48",x"49",x"66",x"c4"),
    73 => (x"a6",x"c8",x"88",x"c1"),
    74 => (x"02",x"99",x"71",x"58"),
    75 => (x"48",x"12",x"87",x"d4"),
    76 => (x"78",x"08",x"d4",x"ff"),
    77 => (x"48",x"49",x"66",x"c4"),
    78 => (x"a6",x"c8",x"88",x"c1"),
    79 => (x"05",x"99",x"71",x"58"),
    80 => (x"4f",x"26",x"87",x"ec"),
    81 => (x"c4",x"4a",x"71",x"1e"),
    82 => (x"c1",x"48",x"49",x"66"),
    83 => (x"58",x"a6",x"c8",x"88"),
    84 => (x"d6",x"02",x"99",x"71"),
    85 => (x"48",x"d4",x"ff",x"87"),
    86 => (x"68",x"78",x"ff",x"c3"),
    87 => (x"49",x"66",x"c4",x"52"),
    88 => (x"c8",x"88",x"c1",x"48"),
    89 => (x"99",x"71",x"58",x"a6"),
    90 => (x"26",x"87",x"ea",x"05"),
    91 => (x"1e",x"73",x"1e",x"4f"),
    92 => (x"c3",x"4b",x"d4",x"ff"),
    93 => (x"4a",x"6b",x"7b",x"ff"),
    94 => (x"6b",x"7b",x"ff",x"c3"),
    95 => (x"72",x"32",x"c8",x"49"),
    96 => (x"7b",x"ff",x"c3",x"b1"),
    97 => (x"31",x"c8",x"4a",x"6b"),
    98 => (x"ff",x"c3",x"b2",x"71"),
    99 => (x"c8",x"49",x"6b",x"7b"),
   100 => (x"71",x"b1",x"72",x"32"),
   101 => (x"26",x"87",x"c4",x"48"),
   102 => (x"26",x"4c",x"26",x"4d"),
   103 => (x"0e",x"4f",x"26",x"4b"),
   104 => (x"5d",x"5c",x"5b",x"5e"),
   105 => (x"ff",x"4a",x"71",x"0e"),
   106 => (x"49",x"72",x"4c",x"d4"),
   107 => (x"71",x"99",x"ff",x"c3"),
   108 => (x"ec",x"e4",x"c2",x"7c"),
   109 => (x"87",x"c8",x"05",x"bf"),
   110 => (x"c9",x"48",x"66",x"d0"),
   111 => (x"58",x"a6",x"d4",x"30"),
   112 => (x"d8",x"49",x"66",x"d0"),
   113 => (x"99",x"ff",x"c3",x"29"),
   114 => (x"66",x"d0",x"7c",x"71"),
   115 => (x"c3",x"29",x"d0",x"49"),
   116 => (x"7c",x"71",x"99",x"ff"),
   117 => (x"c8",x"49",x"66",x"d0"),
   118 => (x"99",x"ff",x"c3",x"29"),
   119 => (x"66",x"d0",x"7c",x"71"),
   120 => (x"99",x"ff",x"c3",x"49"),
   121 => (x"49",x"72",x"7c",x"71"),
   122 => (x"ff",x"c3",x"29",x"d0"),
   123 => (x"6c",x"7c",x"71",x"99"),
   124 => (x"ff",x"f0",x"c9",x"4b"),
   125 => (x"ab",x"ff",x"c3",x"4d"),
   126 => (x"c3",x"87",x"d0",x"05"),
   127 => (x"4b",x"6c",x"7c",x"ff"),
   128 => (x"c6",x"02",x"8d",x"c1"),
   129 => (x"ab",x"ff",x"c3",x"87"),
   130 => (x"73",x"87",x"f0",x"02"),
   131 => (x"87",x"c7",x"fe",x"48"),
   132 => (x"ff",x"49",x"c0",x"1e"),
   133 => (x"ff",x"c3",x"48",x"d4"),
   134 => (x"c3",x"81",x"c1",x"78"),
   135 => (x"04",x"a9",x"b7",x"c8"),
   136 => (x"4f",x"26",x"87",x"f1"),
   137 => (x"e7",x"1e",x"73",x"1e"),
   138 => (x"df",x"f8",x"c4",x"87"),
   139 => (x"c0",x"1e",x"c0",x"4b"),
   140 => (x"f7",x"c1",x"f0",x"ff"),
   141 => (x"87",x"e7",x"fd",x"49"),
   142 => (x"a8",x"c1",x"86",x"c4"),
   143 => (x"87",x"ea",x"c0",x"05"),
   144 => (x"c3",x"48",x"d4",x"ff"),
   145 => (x"c0",x"c1",x"78",x"ff"),
   146 => (x"c0",x"c0",x"c0",x"c0"),
   147 => (x"f0",x"e1",x"c0",x"1e"),
   148 => (x"fd",x"49",x"e9",x"c1"),
   149 => (x"86",x"c4",x"87",x"c9"),
   150 => (x"ca",x"05",x"98",x"70"),
   151 => (x"48",x"d4",x"ff",x"87"),
   152 => (x"c1",x"78",x"ff",x"c3"),
   153 => (x"fe",x"87",x"cb",x"48"),
   154 => (x"8b",x"c1",x"87",x"e6"),
   155 => (x"87",x"fd",x"fe",x"05"),
   156 => (x"e6",x"fc",x"48",x"c0"),
   157 => (x"1e",x"73",x"1e",x"87"),
   158 => (x"c3",x"48",x"d4",x"ff"),
   159 => (x"4b",x"d3",x"78",x"ff"),
   160 => (x"ff",x"c0",x"1e",x"c0"),
   161 => (x"49",x"c1",x"c1",x"f0"),
   162 => (x"c4",x"87",x"d4",x"fc"),
   163 => (x"05",x"98",x"70",x"86"),
   164 => (x"d4",x"ff",x"87",x"ca"),
   165 => (x"78",x"ff",x"c3",x"48"),
   166 => (x"87",x"cb",x"48",x"c1"),
   167 => (x"c1",x"87",x"f1",x"fd"),
   168 => (x"db",x"ff",x"05",x"8b"),
   169 => (x"fb",x"48",x"c0",x"87"),
   170 => (x"5e",x"0e",x"87",x"f1"),
   171 => (x"ff",x"0e",x"5c",x"5b"),
   172 => (x"db",x"fd",x"4c",x"d4"),
   173 => (x"1e",x"ea",x"c6",x"87"),
   174 => (x"c1",x"f0",x"e1",x"c0"),
   175 => (x"de",x"fb",x"49",x"c8"),
   176 => (x"c1",x"86",x"c4",x"87"),
   177 => (x"87",x"c8",x"02",x"a8"),
   178 => (x"c0",x"87",x"ea",x"fe"),
   179 => (x"87",x"e2",x"c1",x"48"),
   180 => (x"70",x"87",x"da",x"fa"),
   181 => (x"ff",x"ff",x"cf",x"49"),
   182 => (x"a9",x"ea",x"c6",x"99"),
   183 => (x"fe",x"87",x"c8",x"02"),
   184 => (x"48",x"c0",x"87",x"d3"),
   185 => (x"c3",x"87",x"cb",x"c1"),
   186 => (x"f1",x"c0",x"7c",x"ff"),
   187 => (x"87",x"f4",x"fc",x"4b"),
   188 => (x"c0",x"02",x"98",x"70"),
   189 => (x"1e",x"c0",x"87",x"eb"),
   190 => (x"c1",x"f0",x"ff",x"c0"),
   191 => (x"de",x"fa",x"49",x"fa"),
   192 => (x"70",x"86",x"c4",x"87"),
   193 => (x"87",x"d9",x"05",x"98"),
   194 => (x"6c",x"7c",x"ff",x"c3"),
   195 => (x"7c",x"ff",x"c3",x"49"),
   196 => (x"c1",x"7c",x"7c",x"7c"),
   197 => (x"c4",x"02",x"99",x"c0"),
   198 => (x"d5",x"48",x"c1",x"87"),
   199 => (x"d1",x"48",x"c0",x"87"),
   200 => (x"05",x"ab",x"c2",x"87"),
   201 => (x"48",x"c0",x"87",x"c4"),
   202 => (x"8b",x"c1",x"87",x"c8"),
   203 => (x"87",x"fd",x"fe",x"05"),
   204 => (x"e4",x"f9",x"48",x"c0"),
   205 => (x"1e",x"73",x"1e",x"87"),
   206 => (x"48",x"ec",x"e4",x"c2"),
   207 => (x"4b",x"c7",x"78",x"c1"),
   208 => (x"c2",x"48",x"d0",x"ff"),
   209 => (x"87",x"c8",x"fb",x"78"),
   210 => (x"c3",x"48",x"d0",x"ff"),
   211 => (x"c0",x"1e",x"c0",x"78"),
   212 => (x"c0",x"c1",x"d0",x"e5"),
   213 => (x"87",x"c7",x"f9",x"49"),
   214 => (x"a8",x"c1",x"86",x"c4"),
   215 => (x"4b",x"87",x"c1",x"05"),
   216 => (x"c5",x"05",x"ab",x"c2"),
   217 => (x"c0",x"48",x"c0",x"87"),
   218 => (x"8b",x"c1",x"87",x"f9"),
   219 => (x"87",x"d0",x"ff",x"05"),
   220 => (x"c2",x"87",x"f7",x"fc"),
   221 => (x"70",x"58",x"f0",x"e4"),
   222 => (x"87",x"cd",x"05",x"98"),
   223 => (x"ff",x"c0",x"1e",x"c1"),
   224 => (x"49",x"d0",x"c1",x"f0"),
   225 => (x"c4",x"87",x"d8",x"f8"),
   226 => (x"48",x"d4",x"ff",x"86"),
   227 => (x"c4",x"78",x"ff",x"c3"),
   228 => (x"e4",x"c2",x"87",x"de"),
   229 => (x"d0",x"ff",x"58",x"f4"),
   230 => (x"ff",x"78",x"c2",x"48"),
   231 => (x"ff",x"c3",x"48",x"d4"),
   232 => (x"f7",x"48",x"c1",x"78"),
   233 => (x"5e",x"0e",x"87",x"f5"),
   234 => (x"0e",x"5d",x"5c",x"5b"),
   235 => (x"ff",x"c3",x"4a",x"71"),
   236 => (x"4c",x"d4",x"ff",x"4d"),
   237 => (x"d0",x"ff",x"7c",x"75"),
   238 => (x"78",x"c3",x"c4",x"48"),
   239 => (x"1e",x"72",x"7c",x"75"),
   240 => (x"c1",x"f0",x"ff",x"c0"),
   241 => (x"d6",x"f7",x"49",x"d8"),
   242 => (x"70",x"86",x"c4",x"87"),
   243 => (x"87",x"c5",x"02",x"98"),
   244 => (x"f0",x"c0",x"48",x"c1"),
   245 => (x"c3",x"7c",x"75",x"87"),
   246 => (x"c0",x"c8",x"7c",x"fe"),
   247 => (x"49",x"66",x"d4",x"1e"),
   248 => (x"c4",x"87",x"fa",x"f4"),
   249 => (x"75",x"7c",x"75",x"86"),
   250 => (x"d8",x"7c",x"75",x"7c"),
   251 => (x"75",x"4b",x"e0",x"da"),
   252 => (x"99",x"49",x"6c",x"7c"),
   253 => (x"c1",x"87",x"c5",x"05"),
   254 => (x"87",x"f3",x"05",x"8b"),
   255 => (x"d0",x"ff",x"7c",x"75"),
   256 => (x"c0",x"78",x"c2",x"48"),
   257 => (x"87",x"cf",x"f6",x"48"),
   258 => (x"5c",x"5b",x"5e",x"0e"),
   259 => (x"4b",x"71",x"0e",x"5d"),
   260 => (x"ee",x"c5",x"4c",x"c0"),
   261 => (x"ff",x"4a",x"df",x"cd"),
   262 => (x"ff",x"c3",x"48",x"d4"),
   263 => (x"c3",x"49",x"68",x"78"),
   264 => (x"c0",x"05",x"a9",x"fe"),
   265 => (x"4d",x"70",x"87",x"fd"),
   266 => (x"cc",x"02",x"9b",x"73"),
   267 => (x"1e",x"66",x"d0",x"87"),
   268 => (x"cf",x"f4",x"49",x"73"),
   269 => (x"d6",x"86",x"c4",x"87"),
   270 => (x"48",x"d0",x"ff",x"87"),
   271 => (x"c3",x"78",x"d1",x"c4"),
   272 => (x"66",x"d0",x"7d",x"ff"),
   273 => (x"d4",x"88",x"c1",x"48"),
   274 => (x"98",x"70",x"58",x"a6"),
   275 => (x"ff",x"87",x"f0",x"05"),
   276 => (x"ff",x"c3",x"48",x"d4"),
   277 => (x"9b",x"73",x"78",x"78"),
   278 => (x"ff",x"87",x"c5",x"05"),
   279 => (x"78",x"d0",x"48",x"d0"),
   280 => (x"c1",x"4c",x"4a",x"c1"),
   281 => (x"ee",x"fe",x"05",x"8a"),
   282 => (x"f4",x"48",x"74",x"87"),
   283 => (x"73",x"1e",x"87",x"e9"),
   284 => (x"c0",x"4a",x"71",x"1e"),
   285 => (x"48",x"d4",x"ff",x"4b"),
   286 => (x"ff",x"78",x"ff",x"c3"),
   287 => (x"c3",x"c4",x"48",x"d0"),
   288 => (x"48",x"d4",x"ff",x"78"),
   289 => (x"72",x"78",x"ff",x"c3"),
   290 => (x"f0",x"ff",x"c0",x"1e"),
   291 => (x"f4",x"49",x"d1",x"c1"),
   292 => (x"86",x"c4",x"87",x"cd"),
   293 => (x"d2",x"05",x"98",x"70"),
   294 => (x"1e",x"c0",x"c8",x"87"),
   295 => (x"fd",x"49",x"66",x"cc"),
   296 => (x"86",x"c4",x"87",x"e6"),
   297 => (x"d0",x"ff",x"4b",x"70"),
   298 => (x"73",x"78",x"c2",x"48"),
   299 => (x"87",x"eb",x"f3",x"48"),
   300 => (x"5c",x"5b",x"5e",x"0e"),
   301 => (x"1e",x"c0",x"0e",x"5d"),
   302 => (x"c1",x"f0",x"ff",x"c0"),
   303 => (x"de",x"f3",x"49",x"c9"),
   304 => (x"c2",x"1e",x"d2",x"87"),
   305 => (x"fc",x"49",x"f4",x"e4"),
   306 => (x"86",x"c8",x"87",x"fe"),
   307 => (x"84",x"c1",x"4c",x"c0"),
   308 => (x"04",x"ac",x"b7",x"d2"),
   309 => (x"e4",x"c2",x"87",x"f8"),
   310 => (x"49",x"bf",x"97",x"f4"),
   311 => (x"c1",x"99",x"c0",x"c3"),
   312 => (x"c0",x"05",x"a9",x"c0"),
   313 => (x"e4",x"c2",x"87",x"e7"),
   314 => (x"49",x"bf",x"97",x"fb"),
   315 => (x"e4",x"c2",x"31",x"d0"),
   316 => (x"4a",x"bf",x"97",x"fc"),
   317 => (x"b1",x"72",x"32",x"c8"),
   318 => (x"97",x"fd",x"e4",x"c2"),
   319 => (x"71",x"b1",x"4a",x"bf"),
   320 => (x"ff",x"ff",x"cf",x"4c"),
   321 => (x"84",x"c1",x"9c",x"ff"),
   322 => (x"e7",x"c1",x"34",x"ca"),
   323 => (x"fd",x"e4",x"c2",x"87"),
   324 => (x"c1",x"49",x"bf",x"97"),
   325 => (x"c2",x"99",x"c6",x"31"),
   326 => (x"bf",x"97",x"fe",x"e4"),
   327 => (x"2a",x"b7",x"c7",x"4a"),
   328 => (x"e4",x"c2",x"b1",x"72"),
   329 => (x"4a",x"bf",x"97",x"f9"),
   330 => (x"c2",x"9d",x"cf",x"4d"),
   331 => (x"bf",x"97",x"fa",x"e4"),
   332 => (x"ca",x"9a",x"c3",x"4a"),
   333 => (x"fb",x"e4",x"c2",x"32"),
   334 => (x"c2",x"4b",x"bf",x"97"),
   335 => (x"c2",x"b2",x"73",x"33"),
   336 => (x"bf",x"97",x"fc",x"e4"),
   337 => (x"9b",x"c0",x"c3",x"4b"),
   338 => (x"73",x"2b",x"b7",x"c6"),
   339 => (x"c1",x"81",x"c2",x"b2"),
   340 => (x"70",x"30",x"71",x"48"),
   341 => (x"75",x"48",x"c1",x"49"),
   342 => (x"72",x"4d",x"70",x"30"),
   343 => (x"71",x"84",x"c1",x"4c"),
   344 => (x"b7",x"c0",x"c8",x"94"),
   345 => (x"87",x"cc",x"06",x"ad"),
   346 => (x"2d",x"b7",x"34",x"c1"),
   347 => (x"ad",x"b7",x"c0",x"c8"),
   348 => (x"87",x"f4",x"ff",x"01"),
   349 => (x"de",x"f0",x"48",x"74"),
   350 => (x"5b",x"5e",x"0e",x"87"),
   351 => (x"f8",x"0e",x"5d",x"5c"),
   352 => (x"da",x"ed",x"c2",x"86"),
   353 => (x"c2",x"78",x"c0",x"48"),
   354 => (x"c0",x"1e",x"d2",x"e5"),
   355 => (x"87",x"de",x"fb",x"49"),
   356 => (x"98",x"70",x"86",x"c4"),
   357 => (x"c0",x"87",x"c5",x"05"),
   358 => (x"87",x"ce",x"c9",x"48"),
   359 => (x"7e",x"c1",x"4d",x"c0"),
   360 => (x"bf",x"c5",x"fa",x"c0"),
   361 => (x"c8",x"e6",x"c2",x"49"),
   362 => (x"4b",x"c8",x"71",x"4a"),
   363 => (x"70",x"87",x"fb",x"ea"),
   364 => (x"87",x"c2",x"05",x"98"),
   365 => (x"fa",x"c0",x"7e",x"c0"),
   366 => (x"c2",x"49",x"bf",x"c1"),
   367 => (x"71",x"4a",x"e4",x"e6"),
   368 => (x"e5",x"ea",x"4b",x"c8"),
   369 => (x"05",x"98",x"70",x"87"),
   370 => (x"7e",x"c0",x"87",x"c2"),
   371 => (x"fd",x"c0",x"02",x"6e"),
   372 => (x"d8",x"ec",x"c2",x"87"),
   373 => (x"ed",x"c2",x"4d",x"bf"),
   374 => (x"7e",x"bf",x"9f",x"d0"),
   375 => (x"ea",x"d6",x"c5",x"48"),
   376 => (x"87",x"c7",x"05",x"a8"),
   377 => (x"bf",x"d8",x"ec",x"c2"),
   378 => (x"6e",x"87",x"ce",x"4d"),
   379 => (x"d5",x"e9",x"ca",x"48"),
   380 => (x"87",x"c5",x"02",x"a8"),
   381 => (x"f1",x"c7",x"48",x"c0"),
   382 => (x"d2",x"e5",x"c2",x"87"),
   383 => (x"f9",x"49",x"75",x"1e"),
   384 => (x"86",x"c4",x"87",x"ec"),
   385 => (x"c5",x"05",x"98",x"70"),
   386 => (x"c7",x"48",x"c0",x"87"),
   387 => (x"fa",x"c0",x"87",x"dc"),
   388 => (x"c2",x"49",x"bf",x"c1"),
   389 => (x"71",x"4a",x"e4",x"e6"),
   390 => (x"cd",x"e9",x"4b",x"c8"),
   391 => (x"05",x"98",x"70",x"87"),
   392 => (x"ed",x"c2",x"87",x"c8"),
   393 => (x"78",x"c1",x"48",x"da"),
   394 => (x"fa",x"c0",x"87",x"da"),
   395 => (x"c2",x"49",x"bf",x"c5"),
   396 => (x"71",x"4a",x"c8",x"e6"),
   397 => (x"f1",x"e8",x"4b",x"c8"),
   398 => (x"02",x"98",x"70",x"87"),
   399 => (x"c0",x"87",x"c5",x"c0"),
   400 => (x"87",x"e6",x"c6",x"48"),
   401 => (x"97",x"d0",x"ed",x"c2"),
   402 => (x"d5",x"c1",x"49",x"bf"),
   403 => (x"cd",x"c0",x"05",x"a9"),
   404 => (x"d1",x"ed",x"c2",x"87"),
   405 => (x"c2",x"49",x"bf",x"97"),
   406 => (x"c0",x"02",x"a9",x"ea"),
   407 => (x"48",x"c0",x"87",x"c5"),
   408 => (x"c2",x"87",x"c7",x"c6"),
   409 => (x"bf",x"97",x"d2",x"e5"),
   410 => (x"e9",x"c3",x"48",x"7e"),
   411 => (x"ce",x"c0",x"02",x"a8"),
   412 => (x"c3",x"48",x"6e",x"87"),
   413 => (x"c0",x"02",x"a8",x"eb"),
   414 => (x"48",x"c0",x"87",x"c5"),
   415 => (x"c2",x"87",x"eb",x"c5"),
   416 => (x"bf",x"97",x"dd",x"e5"),
   417 => (x"c0",x"05",x"99",x"49"),
   418 => (x"e5",x"c2",x"87",x"cc"),
   419 => (x"49",x"bf",x"97",x"de"),
   420 => (x"c0",x"02",x"a9",x"c2"),
   421 => (x"48",x"c0",x"87",x"c5"),
   422 => (x"c2",x"87",x"cf",x"c5"),
   423 => (x"bf",x"97",x"df",x"e5"),
   424 => (x"d6",x"ed",x"c2",x"48"),
   425 => (x"48",x"4c",x"70",x"58"),
   426 => (x"ed",x"c2",x"88",x"c1"),
   427 => (x"e5",x"c2",x"58",x"da"),
   428 => (x"49",x"bf",x"97",x"e0"),
   429 => (x"e5",x"c2",x"81",x"75"),
   430 => (x"4a",x"bf",x"97",x"e1"),
   431 => (x"a1",x"72",x"32",x"c8"),
   432 => (x"e7",x"f1",x"c2",x"7e"),
   433 => (x"c2",x"78",x"6e",x"48"),
   434 => (x"bf",x"97",x"e2",x"e5"),
   435 => (x"58",x"a6",x"c8",x"48"),
   436 => (x"bf",x"da",x"ed",x"c2"),
   437 => (x"87",x"d4",x"c2",x"02"),
   438 => (x"bf",x"c1",x"fa",x"c0"),
   439 => (x"e4",x"e6",x"c2",x"49"),
   440 => (x"4b",x"c8",x"71",x"4a"),
   441 => (x"70",x"87",x"c3",x"e6"),
   442 => (x"c5",x"c0",x"02",x"98"),
   443 => (x"c3",x"48",x"c0",x"87"),
   444 => (x"ed",x"c2",x"87",x"f8"),
   445 => (x"c2",x"4c",x"bf",x"d2"),
   446 => (x"c2",x"5c",x"fb",x"f1"),
   447 => (x"bf",x"97",x"f7",x"e5"),
   448 => (x"c2",x"31",x"c8",x"49"),
   449 => (x"bf",x"97",x"f6",x"e5"),
   450 => (x"c2",x"49",x"a1",x"4a"),
   451 => (x"bf",x"97",x"f8",x"e5"),
   452 => (x"72",x"32",x"d0",x"4a"),
   453 => (x"e5",x"c2",x"49",x"a1"),
   454 => (x"4a",x"bf",x"97",x"f9"),
   455 => (x"a1",x"72",x"32",x"d8"),
   456 => (x"91",x"66",x"c4",x"49"),
   457 => (x"bf",x"e7",x"f1",x"c2"),
   458 => (x"ef",x"f1",x"c2",x"81"),
   459 => (x"ff",x"e5",x"c2",x"59"),
   460 => (x"c8",x"4a",x"bf",x"97"),
   461 => (x"fe",x"e5",x"c2",x"32"),
   462 => (x"a2",x"4b",x"bf",x"97"),
   463 => (x"c0",x"e6",x"c2",x"4a"),
   464 => (x"d0",x"4b",x"bf",x"97"),
   465 => (x"4a",x"a2",x"73",x"33"),
   466 => (x"97",x"c1",x"e6",x"c2"),
   467 => (x"9b",x"cf",x"4b",x"bf"),
   468 => (x"a2",x"73",x"33",x"d8"),
   469 => (x"f3",x"f1",x"c2",x"4a"),
   470 => (x"ef",x"f1",x"c2",x"5a"),
   471 => (x"8a",x"c2",x"4a",x"bf"),
   472 => (x"f1",x"c2",x"92",x"74"),
   473 => (x"a1",x"72",x"48",x"f3"),
   474 => (x"87",x"ca",x"c1",x"78"),
   475 => (x"97",x"e4",x"e5",x"c2"),
   476 => (x"31",x"c8",x"49",x"bf"),
   477 => (x"97",x"e3",x"e5",x"c2"),
   478 => (x"49",x"a1",x"4a",x"bf"),
   479 => (x"59",x"e2",x"ed",x"c2"),
   480 => (x"bf",x"de",x"ed",x"c2"),
   481 => (x"c7",x"31",x"c5",x"49"),
   482 => (x"29",x"c9",x"81",x"ff"),
   483 => (x"59",x"fb",x"f1",x"c2"),
   484 => (x"97",x"e9",x"e5",x"c2"),
   485 => (x"32",x"c8",x"4a",x"bf"),
   486 => (x"97",x"e8",x"e5",x"c2"),
   487 => (x"4a",x"a2",x"4b",x"bf"),
   488 => (x"6e",x"92",x"66",x"c4"),
   489 => (x"f7",x"f1",x"c2",x"82"),
   490 => (x"ef",x"f1",x"c2",x"5a"),
   491 => (x"c2",x"78",x"c0",x"48"),
   492 => (x"72",x"48",x"eb",x"f1"),
   493 => (x"f1",x"c2",x"78",x"a1"),
   494 => (x"f1",x"c2",x"48",x"fb"),
   495 => (x"c2",x"78",x"bf",x"ef"),
   496 => (x"c2",x"48",x"ff",x"f1"),
   497 => (x"78",x"bf",x"f3",x"f1"),
   498 => (x"bf",x"da",x"ed",x"c2"),
   499 => (x"87",x"c9",x"c0",x"02"),
   500 => (x"30",x"c4",x"48",x"74"),
   501 => (x"c9",x"c0",x"7e",x"70"),
   502 => (x"f7",x"f1",x"c2",x"87"),
   503 => (x"30",x"c4",x"48",x"bf"),
   504 => (x"ed",x"c2",x"7e",x"70"),
   505 => (x"78",x"6e",x"48",x"de"),
   506 => (x"8e",x"f8",x"48",x"c1"),
   507 => (x"4c",x"26",x"4d",x"26"),
   508 => (x"4f",x"26",x"4b",x"26"),
   509 => (x"5c",x"5b",x"5e",x"0e"),
   510 => (x"4a",x"71",x"0e",x"5d"),
   511 => (x"bf",x"da",x"ed",x"c2"),
   512 => (x"72",x"87",x"cb",x"02"),
   513 => (x"72",x"2b",x"c7",x"4b"),
   514 => (x"9c",x"ff",x"c1",x"4c"),
   515 => (x"4b",x"72",x"87",x"c9"),
   516 => (x"4c",x"72",x"2b",x"c8"),
   517 => (x"c2",x"9c",x"ff",x"c3"),
   518 => (x"83",x"bf",x"e7",x"f1"),
   519 => (x"bf",x"fd",x"f9",x"c0"),
   520 => (x"87",x"d9",x"02",x"ab"),
   521 => (x"5b",x"c1",x"fa",x"c0"),
   522 => (x"1e",x"d2",x"e5",x"c2"),
   523 => (x"fd",x"f0",x"49",x"73"),
   524 => (x"70",x"86",x"c4",x"87"),
   525 => (x"87",x"c5",x"05",x"98"),
   526 => (x"e6",x"c0",x"48",x"c0"),
   527 => (x"da",x"ed",x"c2",x"87"),
   528 => (x"87",x"d2",x"02",x"bf"),
   529 => (x"91",x"c4",x"49",x"74"),
   530 => (x"81",x"d2",x"e5",x"c2"),
   531 => (x"ff",x"cf",x"4d",x"69"),
   532 => (x"9d",x"ff",x"ff",x"ff"),
   533 => (x"49",x"74",x"87",x"cb"),
   534 => (x"e5",x"c2",x"91",x"c2"),
   535 => (x"69",x"9f",x"81",x"d2"),
   536 => (x"fe",x"48",x"75",x"4d"),
   537 => (x"5e",x"0e",x"87",x"c6"),
   538 => (x"0e",x"5d",x"5c",x"5b"),
   539 => (x"4c",x"71",x"86",x"f4"),
   540 => (x"87",x"c5",x"05",x"9c"),
   541 => (x"f5",x"c3",x"48",x"c0"),
   542 => (x"7e",x"a4",x"c8",x"87"),
   543 => (x"78",x"c0",x"48",x"6e"),
   544 => (x"c7",x"02",x"66",x"dc"),
   545 => (x"97",x"66",x"dc",x"87"),
   546 => (x"87",x"c5",x"05",x"bf"),
   547 => (x"dd",x"c3",x"48",x"c0"),
   548 => (x"c1",x"1e",x"c0",x"87"),
   549 => (x"87",x"c9",x"d0",x"49"),
   550 => (x"a6",x"c8",x"86",x"c4"),
   551 => (x"02",x"66",x"c4",x"58"),
   552 => (x"c2",x"87",x"ff",x"c0"),
   553 => (x"dc",x"4a",x"e2",x"ed"),
   554 => (x"de",x"ff",x"49",x"66"),
   555 => (x"98",x"70",x"87",x"e1"),
   556 => (x"87",x"ee",x"c0",x"02"),
   557 => (x"dc",x"4a",x"66",x"c4"),
   558 => (x"4b",x"cb",x"49",x"66"),
   559 => (x"87",x"c4",x"df",x"ff"),
   560 => (x"dd",x"02",x"98",x"70"),
   561 => (x"c8",x"1e",x"c0",x"87"),
   562 => (x"87",x"c4",x"02",x"66"),
   563 => (x"87",x"c2",x"4d",x"c0"),
   564 => (x"49",x"75",x"4d",x"c1"),
   565 => (x"c4",x"87",x"ca",x"cf"),
   566 => (x"58",x"a6",x"c8",x"86"),
   567 => (x"ff",x"05",x"66",x"c4"),
   568 => (x"66",x"c4",x"87",x"c1"),
   569 => (x"87",x"c4",x"c2",x"02"),
   570 => (x"6e",x"81",x"dc",x"49"),
   571 => (x"c4",x"78",x"69",x"48"),
   572 => (x"81",x"da",x"49",x"66"),
   573 => (x"9f",x"4d",x"a4",x"c4"),
   574 => (x"ed",x"c2",x"7d",x"69"),
   575 => (x"d5",x"02",x"bf",x"da"),
   576 => (x"49",x"66",x"c4",x"87"),
   577 => (x"69",x"9f",x"81",x"d4"),
   578 => (x"ff",x"ff",x"c0",x"49"),
   579 => (x"d0",x"48",x"71",x"99"),
   580 => (x"58",x"a6",x"cc",x"30"),
   581 => (x"a6",x"c8",x"87",x"c5"),
   582 => (x"c8",x"78",x"c0",x"48"),
   583 => (x"6d",x"48",x"49",x"66"),
   584 => (x"c0",x"7d",x"70",x"80"),
   585 => (x"49",x"a4",x"cc",x"7c"),
   586 => (x"a4",x"d0",x"79",x"6d"),
   587 => (x"c4",x"79",x"c0",x"49"),
   588 => (x"78",x"c0",x"48",x"a6"),
   589 => (x"c4",x"4a",x"a4",x"d4"),
   590 => (x"91",x"c8",x"49",x"66"),
   591 => (x"c0",x"49",x"a1",x"72"),
   592 => (x"c4",x"79",x"6d",x"41"),
   593 => (x"80",x"c1",x"48",x"66"),
   594 => (x"c6",x"58",x"a6",x"c8"),
   595 => (x"ff",x"04",x"a8",x"b7"),
   596 => (x"bf",x"6e",x"87",x"e2"),
   597 => (x"72",x"2a",x"c9",x"4a"),
   598 => (x"4a",x"f0",x"c0",x"49"),
   599 => (x"87",x"d8",x"dd",x"ff"),
   600 => (x"c4",x"c1",x"4a",x"70"),
   601 => (x"79",x"72",x"49",x"a4"),
   602 => (x"87",x"c2",x"48",x"c1"),
   603 => (x"8e",x"f4",x"48",x"c0"),
   604 => (x"0e",x"87",x"f9",x"f9"),
   605 => (x"5d",x"5c",x"5b",x"5e"),
   606 => (x"9c",x"4c",x"71",x"0e"),
   607 => (x"87",x"ca",x"c1",x"02"),
   608 => (x"69",x"49",x"a4",x"c8"),
   609 => (x"87",x"c2",x"c1",x"02"),
   610 => (x"6c",x"4a",x"66",x"d0"),
   611 => (x"a6",x"d4",x"82",x"49"),
   612 => (x"4d",x"66",x"d0",x"5a"),
   613 => (x"d6",x"ed",x"c2",x"b9"),
   614 => (x"ba",x"ff",x"4a",x"bf"),
   615 => (x"99",x"71",x"99",x"72"),
   616 => (x"87",x"e4",x"c0",x"02"),
   617 => (x"6b",x"4b",x"a4",x"c4"),
   618 => (x"87",x"c8",x"f9",x"49"),
   619 => (x"ed",x"c2",x"7b",x"70"),
   620 => (x"6c",x"49",x"bf",x"d2"),
   621 => (x"75",x"7c",x"71",x"81"),
   622 => (x"d6",x"ed",x"c2",x"b9"),
   623 => (x"ba",x"ff",x"4a",x"bf"),
   624 => (x"99",x"71",x"99",x"72"),
   625 => (x"87",x"dc",x"ff",x"05"),
   626 => (x"df",x"f8",x"7c",x"75"),
   627 => (x"1e",x"73",x"1e",x"87"),
   628 => (x"02",x"9b",x"4b",x"71"),
   629 => (x"a3",x"c8",x"87",x"c7"),
   630 => (x"c5",x"05",x"69",x"49"),
   631 => (x"c0",x"48",x"c0",x"87"),
   632 => (x"f1",x"c2",x"87",x"f7"),
   633 => (x"c4",x"4a",x"bf",x"eb"),
   634 => (x"49",x"69",x"49",x"a3"),
   635 => (x"ed",x"c2",x"89",x"c2"),
   636 => (x"71",x"91",x"bf",x"d2"),
   637 => (x"ed",x"c2",x"4a",x"a2"),
   638 => (x"6b",x"49",x"bf",x"d6"),
   639 => (x"4a",x"a2",x"71",x"99"),
   640 => (x"5a",x"c1",x"fa",x"c0"),
   641 => (x"72",x"1e",x"66",x"c8"),
   642 => (x"87",x"e2",x"e9",x"49"),
   643 => (x"98",x"70",x"86",x"c4"),
   644 => (x"c0",x"87",x"c4",x"05"),
   645 => (x"c1",x"87",x"c2",x"48"),
   646 => (x"87",x"d4",x"f7",x"48"),
   647 => (x"71",x"1e",x"73",x"1e"),
   648 => (x"c7",x"02",x"9b",x"4b"),
   649 => (x"49",x"a3",x"c8",x"87"),
   650 => (x"87",x"c5",x"05",x"69"),
   651 => (x"f7",x"c0",x"48",x"c0"),
   652 => (x"eb",x"f1",x"c2",x"87"),
   653 => (x"a3",x"c4",x"4a",x"bf"),
   654 => (x"c2",x"49",x"69",x"49"),
   655 => (x"d2",x"ed",x"c2",x"89"),
   656 => (x"a2",x"71",x"91",x"bf"),
   657 => (x"d6",x"ed",x"c2",x"4a"),
   658 => (x"99",x"6b",x"49",x"bf"),
   659 => (x"c0",x"4a",x"a2",x"71"),
   660 => (x"c8",x"5a",x"c1",x"fa"),
   661 => (x"49",x"72",x"1e",x"66"),
   662 => (x"c4",x"87",x"cb",x"e5"),
   663 => (x"05",x"98",x"70",x"86"),
   664 => (x"48",x"c0",x"87",x"c4"),
   665 => (x"48",x"c1",x"87",x"c2"),
   666 => (x"0e",x"87",x"c5",x"f6"),
   667 => (x"5d",x"5c",x"5b",x"5e"),
   668 => (x"71",x"86",x"f8",x"0e"),
   669 => (x"c4",x"7e",x"ff",x"4c"),
   670 => (x"ff",x"c1",x"48",x"a6"),
   671 => (x"ff",x"ff",x"ff",x"ff"),
   672 => (x"d4",x"4b",x"c0",x"78"),
   673 => (x"49",x"73",x"4a",x"a4"),
   674 => (x"a1",x"72",x"91",x"c8"),
   675 => (x"48",x"66",x"d8",x"49"),
   676 => (x"49",x"70",x"88",x"69"),
   677 => (x"ad",x"b7",x"c0",x"4d"),
   678 => (x"c4",x"87",x"cc",x"04"),
   679 => (x"03",x"ad",x"b7",x"66"),
   680 => (x"7e",x"73",x"87",x"c5"),
   681 => (x"c1",x"5d",x"a6",x"c8"),
   682 => (x"ab",x"b7",x"c6",x"83"),
   683 => (x"87",x"d3",x"ff",x"04"),
   684 => (x"8e",x"f8",x"48",x"6e"),
   685 => (x"0e",x"87",x"f5",x"f4"),
   686 => (x"5d",x"5c",x"5b",x"5e"),
   687 => (x"71",x"86",x"f0",x"0e"),
   688 => (x"48",x"a6",x"c4",x"7e"),
   689 => (x"ff",x"ff",x"ff",x"c1"),
   690 => (x"c4",x"78",x"ff",x"ff"),
   691 => (x"c0",x"78",x"ff",x"80"),
   692 => (x"6e",x"4c",x"c0",x"4d"),
   693 => (x"74",x"83",x"d4",x"4b"),
   694 => (x"73",x"92",x"c8",x"4a"),
   695 => (x"49",x"75",x"4a",x"a2"),
   696 => (x"a1",x"73",x"91",x"c8"),
   697 => (x"69",x"48",x"6a",x"49"),
   698 => (x"d0",x"49",x"70",x"88"),
   699 => (x"ad",x"74",x"59",x"a6"),
   700 => (x"cc",x"87",x"cf",x"02"),
   701 => (x"66",x"c4",x"49",x"66"),
   702 => (x"87",x"c6",x"03",x"a9"),
   703 => (x"c8",x"5c",x"a6",x"cc"),
   704 => (x"84",x"c1",x"59",x"a6"),
   705 => (x"04",x"ac",x"b7",x"c6"),
   706 => (x"c1",x"87",x"c8",x"ff"),
   707 => (x"ad",x"b7",x"c6",x"85"),
   708 => (x"87",x"fd",x"fe",x"04"),
   709 => (x"f0",x"48",x"66",x"c8"),
   710 => (x"87",x"d0",x"f3",x"8e"),
   711 => (x"5c",x"5b",x"5e",x"0e"),
   712 => (x"86",x"ec",x"0e",x"5d"),
   713 => (x"e4",x"c0",x"4b",x"71"),
   714 => (x"28",x"c9",x"48",x"66"),
   715 => (x"c2",x"58",x"a6",x"c8"),
   716 => (x"4a",x"bf",x"d6",x"ed"),
   717 => (x"48",x"72",x"ba",x"ff"),
   718 => (x"cc",x"98",x"66",x"c4"),
   719 => (x"9b",x"73",x"58",x"a6"),
   720 => (x"87",x"c2",x"c3",x"02"),
   721 => (x"69",x"49",x"a3",x"c8"),
   722 => (x"87",x"fa",x"c2",x"02"),
   723 => (x"98",x"6b",x"48",x"72"),
   724 => (x"c4",x"58",x"a6",x"d0"),
   725 => (x"7e",x"6c",x"4c",x"a3"),
   726 => (x"cc",x"48",x"66",x"c8"),
   727 => (x"c6",x"05",x"a8",x"66"),
   728 => (x"7b",x"66",x"c4",x"87"),
   729 => (x"c8",x"87",x"cd",x"c2"),
   730 => (x"49",x"73",x"1e",x"66"),
   731 => (x"c4",x"87",x"fc",x"fb"),
   732 => (x"c0",x"4d",x"70",x"86"),
   733 => (x"d0",x"04",x"ad",x"b7"),
   734 => (x"4a",x"a3",x"d4",x"87"),
   735 => (x"91",x"c8",x"49",x"75"),
   736 => (x"21",x"49",x"a1",x"72"),
   737 => (x"c7",x"7c",x"69",x"7b"),
   738 => (x"cc",x"7b",x"c0",x"87"),
   739 => (x"7c",x"69",x"49",x"a3"),
   740 => (x"6b",x"48",x"66",x"c4"),
   741 => (x"58",x"a6",x"c8",x"88"),
   742 => (x"73",x"1e",x"66",x"cc"),
   743 => (x"87",x"cb",x"fb",x"49"),
   744 => (x"4d",x"70",x"86",x"c4"),
   745 => (x"49",x"a3",x"c4",x"c1"),
   746 => (x"69",x"48",x"a6",x"d0"),
   747 => (x"48",x"66",x"cc",x"78"),
   748 => (x"06",x"a8",x"66",x"d0"),
   749 => (x"c0",x"87",x"f2",x"c0"),
   750 => (x"c0",x"04",x"ad",x"b7"),
   751 => (x"a6",x"c8",x"87",x"eb"),
   752 => (x"78",x"a3",x"d4",x"48"),
   753 => (x"91",x"c8",x"49",x"75"),
   754 => (x"cc",x"81",x"66",x"c8"),
   755 => (x"88",x"69",x"48",x"66"),
   756 => (x"66",x"d0",x"49",x"70"),
   757 => (x"87",x"d1",x"06",x"a9"),
   758 => (x"da",x"fb",x"49",x"73"),
   759 => (x"c8",x"49",x"70",x"87"),
   760 => (x"81",x"66",x"c8",x"91"),
   761 => (x"6e",x"41",x"66",x"cc"),
   762 => (x"49",x"66",x"c4",x"79"),
   763 => (x"f6",x"49",x"73",x"1e"),
   764 => (x"86",x"c4",x"87",x"c1"),
   765 => (x"1e",x"d2",x"e5",x"c2"),
   766 => (x"d0",x"f7",x"49",x"73"),
   767 => (x"d0",x"86",x"c4",x"87"),
   768 => (x"e4",x"c0",x"49",x"a3"),
   769 => (x"8e",x"ec",x"79",x"66"),
   770 => (x"1e",x"87",x"e1",x"ef"),
   771 => (x"4b",x"71",x"1e",x"73"),
   772 => (x"e4",x"c0",x"02",x"9b"),
   773 => (x"ff",x"f1",x"c2",x"87"),
   774 => (x"c2",x"4a",x"73",x"5b"),
   775 => (x"d2",x"ed",x"c2",x"8a"),
   776 => (x"c2",x"92",x"49",x"bf"),
   777 => (x"48",x"bf",x"eb",x"f1"),
   778 => (x"f2",x"c2",x"80",x"72"),
   779 => (x"48",x"71",x"58",x"c3"),
   780 => (x"ed",x"c2",x"30",x"c4"),
   781 => (x"ed",x"c0",x"58",x"e2"),
   782 => (x"fb",x"f1",x"c2",x"87"),
   783 => (x"ef",x"f1",x"c2",x"48"),
   784 => (x"f1",x"c2",x"78",x"bf"),
   785 => (x"f1",x"c2",x"48",x"ff"),
   786 => (x"c2",x"78",x"bf",x"f3"),
   787 => (x"02",x"bf",x"da",x"ed"),
   788 => (x"ed",x"c2",x"87",x"c9"),
   789 => (x"c4",x"49",x"bf",x"d2"),
   790 => (x"c2",x"87",x"c7",x"31"),
   791 => (x"49",x"bf",x"f7",x"f1"),
   792 => (x"ed",x"c2",x"31",x"c4"),
   793 => (x"c7",x"ee",x"59",x"e2"),
   794 => (x"5b",x"5e",x"0e",x"87"),
   795 => (x"4a",x"71",x"0e",x"5c"),
   796 => (x"9a",x"72",x"4b",x"c0"),
   797 => (x"87",x"e1",x"c0",x"02"),
   798 => (x"9f",x"49",x"a2",x"da"),
   799 => (x"ed",x"c2",x"4b",x"69"),
   800 => (x"cf",x"02",x"bf",x"da"),
   801 => (x"49",x"a2",x"d4",x"87"),
   802 => (x"4c",x"49",x"69",x"9f"),
   803 => (x"9c",x"ff",x"ff",x"c0"),
   804 => (x"87",x"c2",x"34",x"d0"),
   805 => (x"49",x"74",x"4c",x"c0"),
   806 => (x"fd",x"49",x"73",x"b3"),
   807 => (x"cd",x"ed",x"87",x"ed"),
   808 => (x"5b",x"5e",x"0e",x"87"),
   809 => (x"f4",x"0e",x"5d",x"5c"),
   810 => (x"c0",x"4a",x"71",x"86"),
   811 => (x"02",x"9a",x"72",x"7e"),
   812 => (x"e5",x"c2",x"87",x"d8"),
   813 => (x"78",x"c0",x"48",x"ce"),
   814 => (x"48",x"c6",x"e5",x"c2"),
   815 => (x"bf",x"ff",x"f1",x"c2"),
   816 => (x"ca",x"e5",x"c2",x"78"),
   817 => (x"fb",x"f1",x"c2",x"48"),
   818 => (x"ed",x"c2",x"78",x"bf"),
   819 => (x"50",x"c0",x"48",x"ef"),
   820 => (x"bf",x"de",x"ed",x"c2"),
   821 => (x"ce",x"e5",x"c2",x"49"),
   822 => (x"aa",x"71",x"4a",x"bf"),
   823 => (x"87",x"ca",x"c4",x"03"),
   824 => (x"99",x"cf",x"49",x"72"),
   825 => (x"87",x"ea",x"c0",x"05"),
   826 => (x"48",x"fd",x"f9",x"c0"),
   827 => (x"bf",x"c6",x"e5",x"c2"),
   828 => (x"d2",x"e5",x"c2",x"78"),
   829 => (x"c6",x"e5",x"c2",x"1e"),
   830 => (x"e5",x"c2",x"49",x"bf"),
   831 => (x"a1",x"c1",x"48",x"c6"),
   832 => (x"dd",x"ff",x"71",x"78"),
   833 => (x"86",x"c4",x"87",x"e8"),
   834 => (x"48",x"f9",x"f9",x"c0"),
   835 => (x"78",x"d2",x"e5",x"c2"),
   836 => (x"f9",x"c0",x"87",x"cc"),
   837 => (x"c0",x"48",x"bf",x"f9"),
   838 => (x"f9",x"c0",x"80",x"e0"),
   839 => (x"e5",x"c2",x"58",x"fd"),
   840 => (x"c1",x"48",x"bf",x"ce"),
   841 => (x"d2",x"e5",x"c2",x"80"),
   842 => (x"0e",x"79",x"27",x"58"),
   843 => (x"97",x"bf",x"00",x"00"),
   844 => (x"02",x"9d",x"4d",x"bf"),
   845 => (x"c3",x"87",x"e3",x"c2"),
   846 => (x"c2",x"02",x"ad",x"e5"),
   847 => (x"f9",x"c0",x"87",x"dc"),
   848 => (x"cb",x"4b",x"bf",x"f9"),
   849 => (x"4c",x"11",x"49",x"a3"),
   850 => (x"c1",x"05",x"ac",x"cf"),
   851 => (x"49",x"75",x"87",x"d2"),
   852 => (x"89",x"c1",x"99",x"df"),
   853 => (x"ed",x"c2",x"91",x"cd"),
   854 => (x"a3",x"c1",x"81",x"e2"),
   855 => (x"c3",x"51",x"12",x"4a"),
   856 => (x"51",x"12",x"4a",x"a3"),
   857 => (x"12",x"4a",x"a3",x"c5"),
   858 => (x"4a",x"a3",x"c7",x"51"),
   859 => (x"a3",x"c9",x"51",x"12"),
   860 => (x"ce",x"51",x"12",x"4a"),
   861 => (x"51",x"12",x"4a",x"a3"),
   862 => (x"12",x"4a",x"a3",x"d0"),
   863 => (x"4a",x"a3",x"d2",x"51"),
   864 => (x"a3",x"d4",x"51",x"12"),
   865 => (x"d6",x"51",x"12",x"4a"),
   866 => (x"51",x"12",x"4a",x"a3"),
   867 => (x"12",x"4a",x"a3",x"d8"),
   868 => (x"4a",x"a3",x"dc",x"51"),
   869 => (x"a3",x"de",x"51",x"12"),
   870 => (x"c1",x"51",x"12",x"4a"),
   871 => (x"87",x"fa",x"c0",x"7e"),
   872 => (x"99",x"c8",x"49",x"74"),
   873 => (x"87",x"eb",x"c0",x"05"),
   874 => (x"99",x"d0",x"49",x"74"),
   875 => (x"dc",x"87",x"d1",x"05"),
   876 => (x"cb",x"c0",x"02",x"66"),
   877 => (x"dc",x"49",x"73",x"87"),
   878 => (x"98",x"70",x"0f",x"66"),
   879 => (x"87",x"d3",x"c0",x"02"),
   880 => (x"c6",x"c0",x"05",x"6e"),
   881 => (x"e2",x"ed",x"c2",x"87"),
   882 => (x"c0",x"50",x"c0",x"48"),
   883 => (x"48",x"bf",x"f9",x"f9"),
   884 => (x"c2",x"87",x"e1",x"c2"),
   885 => (x"c0",x"48",x"ef",x"ed"),
   886 => (x"ed",x"c2",x"7e",x"50"),
   887 => (x"c2",x"49",x"bf",x"de"),
   888 => (x"4a",x"bf",x"ce",x"e5"),
   889 => (x"fb",x"04",x"aa",x"71"),
   890 => (x"f1",x"c2",x"87",x"f6"),
   891 => (x"c0",x"05",x"bf",x"ff"),
   892 => (x"ed",x"c2",x"87",x"c8"),
   893 => (x"c1",x"02",x"bf",x"da"),
   894 => (x"e5",x"c2",x"87",x"f8"),
   895 => (x"e7",x"49",x"bf",x"ca"),
   896 => (x"49",x"70",x"87",x"f2"),
   897 => (x"59",x"ce",x"e5",x"c2"),
   898 => (x"c2",x"48",x"a6",x"c4"),
   899 => (x"78",x"bf",x"ca",x"e5"),
   900 => (x"bf",x"da",x"ed",x"c2"),
   901 => (x"87",x"d8",x"c0",x"02"),
   902 => (x"cf",x"49",x"66",x"c4"),
   903 => (x"f8",x"ff",x"ff",x"ff"),
   904 => (x"c0",x"02",x"a9",x"99"),
   905 => (x"4c",x"c0",x"87",x"c5"),
   906 => (x"c1",x"87",x"e1",x"c0"),
   907 => (x"87",x"dc",x"c0",x"4c"),
   908 => (x"cf",x"49",x"66",x"c4"),
   909 => (x"a9",x"99",x"f8",x"ff"),
   910 => (x"87",x"c8",x"c0",x"02"),
   911 => (x"c0",x"48",x"a6",x"c8"),
   912 => (x"87",x"c5",x"c0",x"78"),
   913 => (x"c1",x"48",x"a6",x"c8"),
   914 => (x"4c",x"66",x"c8",x"78"),
   915 => (x"c0",x"05",x"9c",x"74"),
   916 => (x"66",x"c4",x"87",x"e0"),
   917 => (x"c2",x"89",x"c2",x"49"),
   918 => (x"4a",x"bf",x"d2",x"ed"),
   919 => (x"eb",x"f1",x"c2",x"91"),
   920 => (x"e5",x"c2",x"4a",x"bf"),
   921 => (x"a1",x"72",x"48",x"c6"),
   922 => (x"ce",x"e5",x"c2",x"78"),
   923 => (x"f9",x"78",x"c0",x"48"),
   924 => (x"48",x"c0",x"87",x"de"),
   925 => (x"f3",x"e5",x"8e",x"f4"),
   926 => (x"00",x"00",x"00",x"87"),
   927 => (x"ff",x"ff",x"ff",x"00"),
   928 => (x"00",x"0e",x"89",x"ff"),
   929 => (x"00",x"0e",x"92",x"00"),
   930 => (x"54",x"41",x"46",x"00"),
   931 => (x"20",x"20",x"32",x"33"),
   932 => (x"41",x"46",x"00",x"20"),
   933 => (x"20",x"36",x"31",x"54"),
   934 => (x"1e",x"00",x"20",x"20"),
   935 => (x"c3",x"48",x"d4",x"ff"),
   936 => (x"48",x"68",x"78",x"ff"),
   937 => (x"ff",x"1e",x"4f",x"26"),
   938 => (x"ff",x"c3",x"48",x"d4"),
   939 => (x"48",x"d0",x"ff",x"78"),
   940 => (x"ff",x"78",x"e1",x"c0"),
   941 => (x"78",x"d4",x"48",x"d4"),
   942 => (x"48",x"c3",x"f2",x"c2"),
   943 => (x"50",x"bf",x"d4",x"ff"),
   944 => (x"ff",x"1e",x"4f",x"26"),
   945 => (x"e0",x"c0",x"48",x"d0"),
   946 => (x"1e",x"4f",x"26",x"78"),
   947 => (x"70",x"87",x"cc",x"ff"),
   948 => (x"c6",x"02",x"99",x"49"),
   949 => (x"a9",x"fb",x"c0",x"87"),
   950 => (x"71",x"87",x"f1",x"05"),
   951 => (x"0e",x"4f",x"26",x"48"),
   952 => (x"0e",x"5c",x"5b",x"5e"),
   953 => (x"4c",x"c0",x"4b",x"71"),
   954 => (x"70",x"87",x"f0",x"fe"),
   955 => (x"c0",x"02",x"99",x"49"),
   956 => (x"ec",x"c0",x"87",x"f9"),
   957 => (x"f2",x"c0",x"02",x"a9"),
   958 => (x"a9",x"fb",x"c0",x"87"),
   959 => (x"87",x"eb",x"c0",x"02"),
   960 => (x"ac",x"b7",x"66",x"cc"),
   961 => (x"d0",x"87",x"c7",x"03"),
   962 => (x"87",x"c2",x"02",x"66"),
   963 => (x"99",x"71",x"53",x"71"),
   964 => (x"c1",x"87",x"c2",x"02"),
   965 => (x"87",x"c3",x"fe",x"84"),
   966 => (x"02",x"99",x"49",x"70"),
   967 => (x"ec",x"c0",x"87",x"cd"),
   968 => (x"87",x"c7",x"02",x"a9"),
   969 => (x"05",x"a9",x"fb",x"c0"),
   970 => (x"d0",x"87",x"d5",x"ff"),
   971 => (x"87",x"c3",x"02",x"66"),
   972 => (x"c0",x"7b",x"97",x"c0"),
   973 => (x"c4",x"05",x"a9",x"ec"),
   974 => (x"c5",x"4a",x"74",x"87"),
   975 => (x"c0",x"4a",x"74",x"87"),
   976 => (x"48",x"72",x"8a",x"0a"),
   977 => (x"4d",x"26",x"87",x"c2"),
   978 => (x"4b",x"26",x"4c",x"26"),
   979 => (x"fd",x"1e",x"4f",x"26"),
   980 => (x"49",x"70",x"87",x"c9"),
   981 => (x"aa",x"f0",x"c0",x"4a"),
   982 => (x"c0",x"87",x"c9",x"04"),
   983 => (x"c3",x"01",x"aa",x"f9"),
   984 => (x"8a",x"f0",x"c0",x"87"),
   985 => (x"04",x"aa",x"c1",x"c1"),
   986 => (x"da",x"c1",x"87",x"c9"),
   987 => (x"87",x"c3",x"01",x"aa"),
   988 => (x"72",x"8a",x"f7",x"c0"),
   989 => (x"0e",x"4f",x"26",x"48"),
   990 => (x"0e",x"5c",x"5b",x"5e"),
   991 => (x"d4",x"ff",x"4a",x"71"),
   992 => (x"c0",x"49",x"72",x"4c"),
   993 => (x"4b",x"70",x"87",x"e9"),
   994 => (x"87",x"c2",x"02",x"9b"),
   995 => (x"d0",x"ff",x"8b",x"c1"),
   996 => (x"c1",x"78",x"c5",x"48"),
   997 => (x"49",x"73",x"7c",x"d5"),
   998 => (x"ea",x"c1",x"31",x"c6"),
   999 => (x"4a",x"bf",x"97",x"e9"),
  1000 => (x"70",x"b0",x"71",x"48"),
  1001 => (x"48",x"d0",x"ff",x"7c"),
  1002 => (x"48",x"73",x"78",x"c4"),
  1003 => (x"0e",x"87",x"d9",x"fe"),
  1004 => (x"5d",x"5c",x"5b",x"5e"),
  1005 => (x"71",x"86",x"f8",x"0e"),
  1006 => (x"fb",x"7e",x"c0",x"4c"),
  1007 => (x"4b",x"c0",x"87",x"e8"),
  1008 => (x"97",x"dc",x"c1",x"c1"),
  1009 => (x"a9",x"c0",x"49",x"bf"),
  1010 => (x"fb",x"87",x"cf",x"04"),
  1011 => (x"83",x"c1",x"87",x"fd"),
  1012 => (x"97",x"dc",x"c1",x"c1"),
  1013 => (x"06",x"ab",x"49",x"bf"),
  1014 => (x"c1",x"c1",x"87",x"f1"),
  1015 => (x"02",x"bf",x"97",x"dc"),
  1016 => (x"f6",x"fa",x"87",x"cf"),
  1017 => (x"99",x"49",x"70",x"87"),
  1018 => (x"c0",x"87",x"c6",x"02"),
  1019 => (x"f1",x"05",x"a9",x"ec"),
  1020 => (x"fa",x"4b",x"c0",x"87"),
  1021 => (x"4d",x"70",x"87",x"e5"),
  1022 => (x"c8",x"87",x"e0",x"fa"),
  1023 => (x"da",x"fa",x"58",x"a6"),
  1024 => (x"c1",x"4a",x"70",x"87"),
  1025 => (x"49",x"a4",x"c8",x"83"),
  1026 => (x"ad",x"49",x"69",x"97"),
  1027 => (x"c0",x"87",x"c7",x"02"),
  1028 => (x"c0",x"05",x"ad",x"ff"),
  1029 => (x"a4",x"c9",x"87",x"e7"),
  1030 => (x"49",x"69",x"97",x"49"),
  1031 => (x"02",x"a9",x"66",x"c4"),
  1032 => (x"c0",x"48",x"87",x"c7"),
  1033 => (x"d4",x"05",x"a8",x"ff"),
  1034 => (x"49",x"a4",x"ca",x"87"),
  1035 => (x"aa",x"49",x"69",x"97"),
  1036 => (x"c0",x"87",x"c6",x"02"),
  1037 => (x"c4",x"05",x"aa",x"ff"),
  1038 => (x"d0",x"7e",x"c1",x"87"),
  1039 => (x"ad",x"ec",x"c0",x"87"),
  1040 => (x"c0",x"87",x"c6",x"02"),
  1041 => (x"c4",x"05",x"ad",x"fb"),
  1042 => (x"c1",x"4b",x"c0",x"87"),
  1043 => (x"fe",x"02",x"6e",x"7e"),
  1044 => (x"ed",x"f9",x"87",x"e1"),
  1045 => (x"f8",x"48",x"73",x"87"),
  1046 => (x"87",x"ea",x"fb",x"8e"),
  1047 => (x"5b",x"5e",x"0e",x"00"),
  1048 => (x"f8",x"0e",x"5d",x"5c"),
  1049 => (x"ff",x"4d",x"71",x"86"),
  1050 => (x"1e",x"75",x"4b",x"d4"),
  1051 => (x"49",x"c8",x"f2",x"c2"),
  1052 => (x"87",x"f2",x"df",x"ff"),
  1053 => (x"98",x"70",x"86",x"c4"),
  1054 => (x"87",x"cc",x"c4",x"02"),
  1055 => (x"c1",x"48",x"a6",x"c4"),
  1056 => (x"78",x"bf",x"eb",x"ea"),
  1057 => (x"ee",x"fb",x"49",x"75"),
  1058 => (x"48",x"d0",x"ff",x"87"),
  1059 => (x"d6",x"c1",x"78",x"c5"),
  1060 => (x"75",x"4a",x"c0",x"7b"),
  1061 => (x"7b",x"11",x"49",x"a2"),
  1062 => (x"b7",x"cb",x"82",x"c1"),
  1063 => (x"87",x"f3",x"04",x"aa"),
  1064 => (x"ff",x"c3",x"4a",x"cc"),
  1065 => (x"c0",x"82",x"c1",x"7b"),
  1066 => (x"04",x"aa",x"b7",x"e0"),
  1067 => (x"d0",x"ff",x"87",x"f4"),
  1068 => (x"c3",x"78",x"c4",x"48"),
  1069 => (x"78",x"c5",x"7b",x"ff"),
  1070 => (x"c1",x"7b",x"d3",x"c1"),
  1071 => (x"66",x"78",x"c4",x"7b"),
  1072 => (x"a8",x"b7",x"c0",x"48"),
  1073 => (x"87",x"f0",x"c2",x"06"),
  1074 => (x"bf",x"d0",x"f2",x"c2"),
  1075 => (x"48",x"66",x"c4",x"4c"),
  1076 => (x"a6",x"c8",x"88",x"74"),
  1077 => (x"02",x"9c",x"74",x"58"),
  1078 => (x"c2",x"87",x"f9",x"c1"),
  1079 => (x"c8",x"7e",x"d2",x"e5"),
  1080 => (x"c0",x"8c",x"4d",x"c0"),
  1081 => (x"c6",x"03",x"ac",x"b7"),
  1082 => (x"a4",x"c0",x"c8",x"87"),
  1083 => (x"c2",x"4c",x"c0",x"4d"),
  1084 => (x"bf",x"97",x"c3",x"f2"),
  1085 => (x"02",x"99",x"d0",x"49"),
  1086 => (x"1e",x"c0",x"87",x"d1"),
  1087 => (x"49",x"c8",x"f2",x"c2"),
  1088 => (x"c4",x"87",x"ca",x"e3"),
  1089 => (x"4a",x"49",x"70",x"86"),
  1090 => (x"c2",x"87",x"ee",x"c0"),
  1091 => (x"c2",x"1e",x"d2",x"e5"),
  1092 => (x"e2",x"49",x"c8",x"f2"),
  1093 => (x"86",x"c4",x"87",x"f7"),
  1094 => (x"ff",x"4a",x"49",x"70"),
  1095 => (x"c5",x"c8",x"48",x"d0"),
  1096 => (x"7b",x"d4",x"c1",x"78"),
  1097 => (x"7b",x"bf",x"97",x"6e"),
  1098 => (x"80",x"c1",x"48",x"6e"),
  1099 => (x"8d",x"c1",x"7e",x"70"),
  1100 => (x"87",x"f0",x"ff",x"05"),
  1101 => (x"c4",x"48",x"d0",x"ff"),
  1102 => (x"05",x"9a",x"72",x"78"),
  1103 => (x"48",x"c0",x"87",x"c5"),
  1104 => (x"c1",x"87",x"c7",x"c1"),
  1105 => (x"c8",x"f2",x"c2",x"1e"),
  1106 => (x"87",x"e7",x"e0",x"49"),
  1107 => (x"9c",x"74",x"86",x"c4"),
  1108 => (x"87",x"c7",x"fe",x"05"),
  1109 => (x"c0",x"48",x"66",x"c4"),
  1110 => (x"d1",x"06",x"a8",x"b7"),
  1111 => (x"c8",x"f2",x"c2",x"87"),
  1112 => (x"d0",x"78",x"c0",x"48"),
  1113 => (x"f4",x"78",x"c0",x"80"),
  1114 => (x"d4",x"f2",x"c2",x"80"),
  1115 => (x"66",x"c4",x"78",x"bf"),
  1116 => (x"a8",x"b7",x"c0",x"48"),
  1117 => (x"87",x"d0",x"fd",x"01"),
  1118 => (x"c5",x"48",x"d0",x"ff"),
  1119 => (x"7b",x"d3",x"c1",x"78"),
  1120 => (x"78",x"c4",x"7b",x"c0"),
  1121 => (x"87",x"c2",x"48",x"c1"),
  1122 => (x"8e",x"f8",x"48",x"c0"),
  1123 => (x"4c",x"26",x"4d",x"26"),
  1124 => (x"4f",x"26",x"4b",x"26"),
  1125 => (x"5c",x"5b",x"5e",x"0e"),
  1126 => (x"71",x"1e",x"0e",x"5d"),
  1127 => (x"4d",x"4c",x"c0",x"4b"),
  1128 => (x"e8",x"c0",x"04",x"ab"),
  1129 => (x"ef",x"fe",x"c0",x"87"),
  1130 => (x"02",x"9d",x"75",x"1e"),
  1131 => (x"4a",x"c0",x"87",x"c4"),
  1132 => (x"4a",x"c1",x"87",x"c2"),
  1133 => (x"e8",x"eb",x"49",x"72"),
  1134 => (x"70",x"86",x"c4",x"87"),
  1135 => (x"6e",x"84",x"c1",x"7e"),
  1136 => (x"73",x"87",x"c2",x"05"),
  1137 => (x"73",x"85",x"c1",x"4c"),
  1138 => (x"d8",x"ff",x"06",x"ac"),
  1139 => (x"26",x"48",x"6e",x"87"),
  1140 => (x"0e",x"87",x"f9",x"fe"),
  1141 => (x"0e",x"5c",x"5b",x"5e"),
  1142 => (x"66",x"cc",x"4b",x"71"),
  1143 => (x"4c",x"87",x"d8",x"02"),
  1144 => (x"02",x"8c",x"f0",x"c0"),
  1145 => (x"4a",x"74",x"87",x"d8"),
  1146 => (x"d1",x"02",x"8a",x"c1"),
  1147 => (x"cd",x"02",x"8a",x"87"),
  1148 => (x"c9",x"02",x"8a",x"87"),
  1149 => (x"73",x"87",x"d9",x"87"),
  1150 => (x"87",x"e1",x"f9",x"49"),
  1151 => (x"1e",x"74",x"87",x"d2"),
  1152 => (x"d8",x"c1",x"49",x"c0"),
  1153 => (x"1e",x"74",x"87",x"fb"),
  1154 => (x"d8",x"c1",x"49",x"73"),
  1155 => (x"86",x"c8",x"87",x"f3"),
  1156 => (x"0e",x"87",x"fb",x"fd"),
  1157 => (x"5d",x"5c",x"5b",x"5e"),
  1158 => (x"4c",x"71",x"1e",x"0e"),
  1159 => (x"c2",x"91",x"de",x"49"),
  1160 => (x"71",x"4d",x"e4",x"f3"),
  1161 => (x"02",x"6d",x"97",x"85"),
  1162 => (x"c2",x"87",x"dc",x"c1"),
  1163 => (x"4a",x"bf",x"d0",x"f3"),
  1164 => (x"49",x"72",x"82",x"74"),
  1165 => (x"70",x"87",x"dd",x"fd"),
  1166 => (x"c0",x"02",x"6e",x"7e"),
  1167 => (x"f3",x"c2",x"87",x"f2"),
  1168 => (x"4a",x"6e",x"4b",x"d8"),
  1169 => (x"f9",x"fe",x"49",x"cb"),
  1170 => (x"4b",x"74",x"87",x"de"),
  1171 => (x"ea",x"c1",x"93",x"cb"),
  1172 => (x"83",x"c4",x"83",x"fd"),
  1173 => (x"7b",x"cb",x"ca",x"c1"),
  1174 => (x"c1",x"c1",x"49",x"74"),
  1175 => (x"7b",x"75",x"87",x"f0"),
  1176 => (x"97",x"ea",x"ea",x"c1"),
  1177 => (x"c2",x"1e",x"49",x"bf"),
  1178 => (x"fd",x"49",x"d8",x"f3"),
  1179 => (x"86",x"c4",x"87",x"e5"),
  1180 => (x"c1",x"c1",x"49",x"74"),
  1181 => (x"49",x"c0",x"87",x"d8"),
  1182 => (x"87",x"f7",x"c2",x"c1"),
  1183 => (x"48",x"c4",x"f2",x"c2"),
  1184 => (x"49",x"c1",x"78",x"c0"),
  1185 => (x"26",x"87",x"da",x"dd"),
  1186 => (x"4c",x"87",x"c1",x"fc"),
  1187 => (x"69",x"64",x"61",x"6f"),
  1188 => (x"2e",x"2e",x"67",x"6e"),
  1189 => (x"5e",x"0e",x"00",x"2e"),
  1190 => (x"71",x"0e",x"5c",x"5b"),
  1191 => (x"f3",x"c2",x"4a",x"4b"),
  1192 => (x"72",x"82",x"bf",x"d0"),
  1193 => (x"87",x"ec",x"fb",x"49"),
  1194 => (x"02",x"9c",x"4c",x"70"),
  1195 => (x"e6",x"49",x"87",x"c4"),
  1196 => (x"f3",x"c2",x"87",x"f7"),
  1197 => (x"78",x"c0",x"48",x"d0"),
  1198 => (x"e4",x"dc",x"49",x"c1"),
  1199 => (x"87",x"ce",x"fb",x"87"),
  1200 => (x"5c",x"5b",x"5e",x"0e"),
  1201 => (x"86",x"f4",x"0e",x"5d"),
  1202 => (x"4d",x"d2",x"e5",x"c2"),
  1203 => (x"a6",x"c4",x"4c",x"c0"),
  1204 => (x"c2",x"78",x"c0",x"48"),
  1205 => (x"49",x"bf",x"d0",x"f3"),
  1206 => (x"c1",x"06",x"a9",x"c0"),
  1207 => (x"e5",x"c2",x"87",x"c1"),
  1208 => (x"02",x"98",x"48",x"d2"),
  1209 => (x"c0",x"87",x"f8",x"c0"),
  1210 => (x"c8",x"1e",x"ef",x"fe"),
  1211 => (x"87",x"c7",x"02",x"66"),
  1212 => (x"c0",x"48",x"a6",x"c4"),
  1213 => (x"c4",x"87",x"c5",x"78"),
  1214 => (x"78",x"c1",x"48",x"a6"),
  1215 => (x"e6",x"49",x"66",x"c4"),
  1216 => (x"86",x"c4",x"87",x"df"),
  1217 => (x"84",x"c1",x"4d",x"70"),
  1218 => (x"c1",x"48",x"66",x"c4"),
  1219 => (x"58",x"a6",x"c8",x"80"),
  1220 => (x"bf",x"d0",x"f3",x"c2"),
  1221 => (x"c6",x"03",x"ac",x"49"),
  1222 => (x"05",x"9d",x"75",x"87"),
  1223 => (x"c0",x"87",x"c8",x"ff"),
  1224 => (x"02",x"9d",x"75",x"4c"),
  1225 => (x"c0",x"87",x"e0",x"c3"),
  1226 => (x"c8",x"1e",x"ef",x"fe"),
  1227 => (x"87",x"c7",x"02",x"66"),
  1228 => (x"c0",x"48",x"a6",x"cc"),
  1229 => (x"cc",x"87",x"c5",x"78"),
  1230 => (x"78",x"c1",x"48",x"a6"),
  1231 => (x"e5",x"49",x"66",x"cc"),
  1232 => (x"86",x"c4",x"87",x"df"),
  1233 => (x"02",x"6e",x"7e",x"70"),
  1234 => (x"6e",x"87",x"e9",x"c2"),
  1235 => (x"97",x"81",x"cb",x"49"),
  1236 => (x"99",x"d0",x"49",x"69"),
  1237 => (x"87",x"d6",x"c1",x"02"),
  1238 => (x"4a",x"d6",x"ca",x"c1"),
  1239 => (x"91",x"cb",x"49",x"74"),
  1240 => (x"81",x"fd",x"ea",x"c1"),
  1241 => (x"81",x"c8",x"79",x"72"),
  1242 => (x"74",x"51",x"ff",x"c3"),
  1243 => (x"c2",x"91",x"de",x"49"),
  1244 => (x"71",x"4d",x"e4",x"f3"),
  1245 => (x"97",x"c1",x"c2",x"85"),
  1246 => (x"49",x"a5",x"c1",x"7d"),
  1247 => (x"c2",x"51",x"e0",x"c0"),
  1248 => (x"bf",x"97",x"e2",x"ed"),
  1249 => (x"c1",x"87",x"d2",x"02"),
  1250 => (x"4b",x"a5",x"c2",x"84"),
  1251 => (x"4a",x"e2",x"ed",x"c2"),
  1252 => (x"f4",x"fe",x"49",x"db"),
  1253 => (x"db",x"c1",x"87",x"d2"),
  1254 => (x"49",x"a5",x"cd",x"87"),
  1255 => (x"84",x"c1",x"51",x"c0"),
  1256 => (x"6e",x"4b",x"a5",x"c2"),
  1257 => (x"fe",x"49",x"cb",x"4a"),
  1258 => (x"c1",x"87",x"fd",x"f3"),
  1259 => (x"c8",x"c1",x"87",x"c6"),
  1260 => (x"49",x"74",x"4a",x"d3"),
  1261 => (x"ea",x"c1",x"91",x"cb"),
  1262 => (x"79",x"72",x"81",x"fd"),
  1263 => (x"97",x"e2",x"ed",x"c2"),
  1264 => (x"87",x"d8",x"02",x"bf"),
  1265 => (x"91",x"de",x"49",x"74"),
  1266 => (x"f3",x"c2",x"84",x"c1"),
  1267 => (x"83",x"71",x"4b",x"e4"),
  1268 => (x"4a",x"e2",x"ed",x"c2"),
  1269 => (x"f3",x"fe",x"49",x"dd"),
  1270 => (x"87",x"d8",x"87",x"ce"),
  1271 => (x"93",x"de",x"4b",x"74"),
  1272 => (x"83",x"e4",x"f3",x"c2"),
  1273 => (x"c0",x"49",x"a3",x"cb"),
  1274 => (x"73",x"84",x"c1",x"51"),
  1275 => (x"49",x"cb",x"4a",x"6e"),
  1276 => (x"87",x"f4",x"f2",x"fe"),
  1277 => (x"c1",x"48",x"66",x"c4"),
  1278 => (x"58",x"a6",x"c8",x"80"),
  1279 => (x"c0",x"03",x"ac",x"c7"),
  1280 => (x"05",x"6e",x"87",x"c5"),
  1281 => (x"74",x"87",x"e0",x"fc"),
  1282 => (x"f5",x"8e",x"f4",x"48"),
  1283 => (x"73",x"1e",x"87",x"fe"),
  1284 => (x"49",x"4b",x"71",x"1e"),
  1285 => (x"ea",x"c1",x"91",x"cb"),
  1286 => (x"a1",x"c8",x"81",x"fd"),
  1287 => (x"e9",x"ea",x"c1",x"4a"),
  1288 => (x"c9",x"50",x"12",x"48"),
  1289 => (x"c1",x"c1",x"4a",x"a1"),
  1290 => (x"50",x"12",x"48",x"dc"),
  1291 => (x"ea",x"c1",x"81",x"ca"),
  1292 => (x"50",x"11",x"48",x"ea"),
  1293 => (x"97",x"ea",x"ea",x"c1"),
  1294 => (x"c0",x"1e",x"49",x"bf"),
  1295 => (x"87",x"d3",x"f6",x"49"),
  1296 => (x"48",x"c4",x"f2",x"c2"),
  1297 => (x"49",x"c1",x"78",x"de"),
  1298 => (x"26",x"87",x"d6",x"d6"),
  1299 => (x"1e",x"87",x"c1",x"f5"),
  1300 => (x"cb",x"49",x"4a",x"71"),
  1301 => (x"fd",x"ea",x"c1",x"91"),
  1302 => (x"11",x"81",x"c8",x"81"),
  1303 => (x"c8",x"f2",x"c2",x"48"),
  1304 => (x"d0",x"f3",x"c2",x"58"),
  1305 => (x"c1",x"78",x"c0",x"48"),
  1306 => (x"87",x"f5",x"d5",x"49"),
  1307 => (x"c0",x"1e",x"4f",x"26"),
  1308 => (x"fe",x"fa",x"c0",x"49"),
  1309 => (x"1e",x"4f",x"26",x"87"),
  1310 => (x"d2",x"02",x"99",x"71"),
  1311 => (x"d2",x"ec",x"c1",x"87"),
  1312 => (x"f7",x"50",x"c0",x"48"),
  1313 => (x"cf",x"d1",x"c1",x"80"),
  1314 => (x"f6",x"ea",x"c1",x"40"),
  1315 => (x"c1",x"87",x"ce",x"78"),
  1316 => (x"c1",x"48",x"ce",x"ec"),
  1317 => (x"fc",x"78",x"ef",x"ea"),
  1318 => (x"ee",x"d1",x"c1",x"80"),
  1319 => (x"0e",x"4f",x"26",x"78"),
  1320 => (x"0e",x"5c",x"5b",x"5e"),
  1321 => (x"cb",x"4a",x"4c",x"71"),
  1322 => (x"fd",x"ea",x"c1",x"92"),
  1323 => (x"49",x"a2",x"c8",x"82"),
  1324 => (x"97",x"4b",x"a2",x"c9"),
  1325 => (x"97",x"1e",x"4b",x"6b"),
  1326 => (x"ca",x"1e",x"49",x"69"),
  1327 => (x"c0",x"49",x"12",x"82"),
  1328 => (x"c0",x"87",x"f9",x"e5"),
  1329 => (x"87",x"d9",x"d4",x"49"),
  1330 => (x"f8",x"c0",x"49",x"74"),
  1331 => (x"8e",x"f8",x"87",x"c0"),
  1332 => (x"1e",x"87",x"fb",x"f2"),
  1333 => (x"4b",x"71",x"1e",x"73"),
  1334 => (x"87",x"c3",x"ff",x"49"),
  1335 => (x"fe",x"fe",x"49",x"73"),
  1336 => (x"87",x"ec",x"f2",x"87"),
  1337 => (x"71",x"1e",x"73",x"1e"),
  1338 => (x"4a",x"a3",x"c6",x"4b"),
  1339 => (x"c1",x"87",x"db",x"02"),
  1340 => (x"87",x"d6",x"02",x"8a"),
  1341 => (x"da",x"c1",x"02",x"8a"),
  1342 => (x"c0",x"02",x"8a",x"87"),
  1343 => (x"02",x"8a",x"87",x"fc"),
  1344 => (x"8a",x"87",x"e1",x"c0"),
  1345 => (x"c1",x"87",x"cb",x"02"),
  1346 => (x"49",x"c7",x"87",x"db"),
  1347 => (x"c1",x"87",x"c0",x"fd"),
  1348 => (x"f3",x"c2",x"87",x"de"),
  1349 => (x"c1",x"02",x"bf",x"d0"),
  1350 => (x"c1",x"48",x"87",x"cb"),
  1351 => (x"d4",x"f3",x"c2",x"88"),
  1352 => (x"87",x"c1",x"c1",x"58"),
  1353 => (x"bf",x"d4",x"f3",x"c2"),
  1354 => (x"87",x"f9",x"c0",x"02"),
  1355 => (x"bf",x"d0",x"f3",x"c2"),
  1356 => (x"c2",x"80",x"c1",x"48"),
  1357 => (x"c0",x"58",x"d4",x"f3"),
  1358 => (x"f3",x"c2",x"87",x"eb"),
  1359 => (x"c6",x"49",x"bf",x"d0"),
  1360 => (x"d4",x"f3",x"c2",x"89"),
  1361 => (x"a9",x"b7",x"c0",x"59"),
  1362 => (x"c2",x"87",x"da",x"03"),
  1363 => (x"c0",x"48",x"d0",x"f3"),
  1364 => (x"c2",x"87",x"d2",x"78"),
  1365 => (x"02",x"bf",x"d4",x"f3"),
  1366 => (x"f3",x"c2",x"87",x"cb"),
  1367 => (x"c6",x"48",x"bf",x"d0"),
  1368 => (x"d4",x"f3",x"c2",x"80"),
  1369 => (x"d1",x"49",x"c0",x"58"),
  1370 => (x"49",x"73",x"87",x"f7"),
  1371 => (x"87",x"de",x"f5",x"c0"),
  1372 => (x"0e",x"87",x"dd",x"f0"),
  1373 => (x"5d",x"5c",x"5b",x"5e"),
  1374 => (x"86",x"d0",x"ff",x"0e"),
  1375 => (x"c8",x"59",x"a6",x"dc"),
  1376 => (x"78",x"c0",x"48",x"a6"),
  1377 => (x"c4",x"c1",x"80",x"c4"),
  1378 => (x"80",x"c4",x"78",x"66"),
  1379 => (x"80",x"c4",x"78",x"c1"),
  1380 => (x"f3",x"c2",x"78",x"c1"),
  1381 => (x"78",x"c1",x"48",x"d4"),
  1382 => (x"bf",x"c4",x"f2",x"c2"),
  1383 => (x"05",x"a8",x"de",x"48"),
  1384 => (x"db",x"f4",x"87",x"cb"),
  1385 => (x"cc",x"49",x"70",x"87"),
  1386 => (x"f3",x"cf",x"59",x"a6"),
  1387 => (x"87",x"f6",x"e3",x"87"),
  1388 => (x"e3",x"87",x"d8",x"e4"),
  1389 => (x"4c",x"70",x"87",x"e5"),
  1390 => (x"02",x"ac",x"fb",x"c0"),
  1391 => (x"d8",x"87",x"fb",x"c1"),
  1392 => (x"ed",x"c1",x"05",x"66"),
  1393 => (x"66",x"c0",x"c1",x"87"),
  1394 => (x"6a",x"82",x"c4",x"4a"),
  1395 => (x"c1",x"1e",x"72",x"7e"),
  1396 => (x"c4",x"48",x"d5",x"e7"),
  1397 => (x"a1",x"c8",x"49",x"66"),
  1398 => (x"71",x"41",x"20",x"4a"),
  1399 => (x"87",x"f9",x"05",x"aa"),
  1400 => (x"4a",x"26",x"51",x"10"),
  1401 => (x"48",x"66",x"c0",x"c1"),
  1402 => (x"78",x"ce",x"d0",x"c1"),
  1403 => (x"81",x"c7",x"49",x"6a"),
  1404 => (x"c0",x"c1",x"51",x"74"),
  1405 => (x"81",x"c8",x"49",x"66"),
  1406 => (x"c0",x"c1",x"51",x"c1"),
  1407 => (x"81",x"c9",x"49",x"66"),
  1408 => (x"c0",x"c1",x"51",x"c0"),
  1409 => (x"81",x"ca",x"49",x"66"),
  1410 => (x"1e",x"c1",x"51",x"c0"),
  1411 => (x"49",x"6a",x"1e",x"d8"),
  1412 => (x"ca",x"e3",x"81",x"c8"),
  1413 => (x"c1",x"86",x"c8",x"87"),
  1414 => (x"c0",x"48",x"66",x"c4"),
  1415 => (x"87",x"c7",x"01",x"a8"),
  1416 => (x"c1",x"48",x"a6",x"c8"),
  1417 => (x"c1",x"87",x"ce",x"78"),
  1418 => (x"c1",x"48",x"66",x"c4"),
  1419 => (x"58",x"a6",x"d0",x"88"),
  1420 => (x"d6",x"e2",x"87",x"c3"),
  1421 => (x"48",x"a6",x"d0",x"87"),
  1422 => (x"9c",x"74",x"78",x"c2"),
  1423 => (x"87",x"dc",x"cd",x"02"),
  1424 => (x"c1",x"48",x"66",x"c8"),
  1425 => (x"03",x"a8",x"66",x"c8"),
  1426 => (x"dc",x"87",x"d1",x"cd"),
  1427 => (x"78",x"c0",x"48",x"a6"),
  1428 => (x"78",x"c0",x"80",x"e8"),
  1429 => (x"70",x"87",x"c4",x"e1"),
  1430 => (x"ac",x"d0",x"c1",x"4c"),
  1431 => (x"87",x"d8",x"c2",x"05"),
  1432 => (x"e3",x"7e",x"66",x"c4"),
  1433 => (x"49",x"70",x"87",x"e8"),
  1434 => (x"e0",x"59",x"a6",x"c8"),
  1435 => (x"4c",x"70",x"87",x"ed"),
  1436 => (x"05",x"ac",x"ec",x"c0"),
  1437 => (x"c8",x"87",x"ec",x"c1"),
  1438 => (x"91",x"cb",x"49",x"66"),
  1439 => (x"81",x"66",x"c0",x"c1"),
  1440 => (x"6a",x"4a",x"a1",x"c4"),
  1441 => (x"4a",x"a1",x"c8",x"4d"),
  1442 => (x"c1",x"52",x"66",x"c4"),
  1443 => (x"e0",x"79",x"cf",x"d1"),
  1444 => (x"4c",x"70",x"87",x"c9"),
  1445 => (x"87",x"d9",x"02",x"9c"),
  1446 => (x"02",x"ac",x"fb",x"c0"),
  1447 => (x"55",x"74",x"87",x"d3"),
  1448 => (x"87",x"f7",x"df",x"ff"),
  1449 => (x"02",x"9c",x"4c",x"70"),
  1450 => (x"fb",x"c0",x"87",x"c7"),
  1451 => (x"ed",x"ff",x"05",x"ac"),
  1452 => (x"55",x"e0",x"c0",x"87"),
  1453 => (x"c0",x"55",x"c1",x"c2"),
  1454 => (x"66",x"d8",x"7d",x"97"),
  1455 => (x"05",x"a9",x"6e",x"49"),
  1456 => (x"66",x"c8",x"87",x"db"),
  1457 => (x"a8",x"66",x"cc",x"48"),
  1458 => (x"c8",x"87",x"ca",x"04"),
  1459 => (x"80",x"c1",x"48",x"66"),
  1460 => (x"c8",x"58",x"a6",x"cc"),
  1461 => (x"48",x"66",x"cc",x"87"),
  1462 => (x"a6",x"d0",x"88",x"c1"),
  1463 => (x"fa",x"de",x"ff",x"58"),
  1464 => (x"c1",x"4c",x"70",x"87"),
  1465 => (x"c8",x"05",x"ac",x"d0"),
  1466 => (x"48",x"66",x"d4",x"87"),
  1467 => (x"a6",x"d8",x"80",x"c1"),
  1468 => (x"ac",x"d0",x"c1",x"58"),
  1469 => (x"87",x"e8",x"fd",x"02"),
  1470 => (x"48",x"a6",x"e0",x"c0"),
  1471 => (x"c4",x"78",x"66",x"d8"),
  1472 => (x"e0",x"c0",x"48",x"66"),
  1473 => (x"c9",x"05",x"a8",x"66"),
  1474 => (x"e4",x"c0",x"87",x"e4"),
  1475 => (x"78",x"c0",x"48",x"a6"),
  1476 => (x"78",x"c0",x"80",x"c4"),
  1477 => (x"fb",x"c0",x"48",x"74"),
  1478 => (x"6e",x"7e",x"70",x"88"),
  1479 => (x"87",x"e7",x"c8",x"02"),
  1480 => (x"88",x"cb",x"48",x"6e"),
  1481 => (x"02",x"6e",x"7e",x"70"),
  1482 => (x"6e",x"87",x"cd",x"c1"),
  1483 => (x"70",x"88",x"c9",x"48"),
  1484 => (x"c3",x"02",x"6e",x"7e"),
  1485 => (x"48",x"6e",x"87",x"e9"),
  1486 => (x"7e",x"70",x"88",x"c4"),
  1487 => (x"87",x"ce",x"02",x"6e"),
  1488 => (x"88",x"c1",x"48",x"6e"),
  1489 => (x"02",x"6e",x"7e",x"70"),
  1490 => (x"c7",x"87",x"d4",x"c3"),
  1491 => (x"a6",x"dc",x"87",x"f3"),
  1492 => (x"78",x"f0",x"c0",x"48"),
  1493 => (x"87",x"c3",x"dd",x"ff"),
  1494 => (x"ec",x"c0",x"4c",x"70"),
  1495 => (x"c4",x"c0",x"02",x"ac"),
  1496 => (x"a6",x"e0",x"c0",x"87"),
  1497 => (x"ac",x"ec",x"c0",x"5c"),
  1498 => (x"ff",x"87",x"cd",x"02"),
  1499 => (x"70",x"87",x"ec",x"dc"),
  1500 => (x"ac",x"ec",x"c0",x"4c"),
  1501 => (x"87",x"f3",x"ff",x"05"),
  1502 => (x"02",x"ac",x"ec",x"c0"),
  1503 => (x"ff",x"87",x"c4",x"c0"),
  1504 => (x"c0",x"87",x"d8",x"dc"),
  1505 => (x"d0",x"1e",x"ca",x"1e"),
  1506 => (x"91",x"cb",x"49",x"66"),
  1507 => (x"48",x"66",x"c8",x"c1"),
  1508 => (x"a6",x"cc",x"80",x"71"),
  1509 => (x"48",x"66",x"c8",x"58"),
  1510 => (x"a6",x"d0",x"80",x"c4"),
  1511 => (x"bf",x"66",x"cc",x"58"),
  1512 => (x"fa",x"dc",x"ff",x"49"),
  1513 => (x"de",x"1e",x"c1",x"87"),
  1514 => (x"bf",x"66",x"d4",x"1e"),
  1515 => (x"ee",x"dc",x"ff",x"49"),
  1516 => (x"70",x"86",x"d0",x"87"),
  1517 => (x"89",x"09",x"c0",x"49"),
  1518 => (x"59",x"a6",x"ec",x"c0"),
  1519 => (x"48",x"66",x"e8",x"c0"),
  1520 => (x"c0",x"06",x"a8",x"c0"),
  1521 => (x"e8",x"c0",x"87",x"ee"),
  1522 => (x"a8",x"dd",x"48",x"66"),
  1523 => (x"87",x"e4",x"c0",x"03"),
  1524 => (x"49",x"bf",x"66",x"c4"),
  1525 => (x"81",x"66",x"e8",x"c0"),
  1526 => (x"c0",x"51",x"e0",x"c0"),
  1527 => (x"c1",x"49",x"66",x"e8"),
  1528 => (x"bf",x"66",x"c4",x"81"),
  1529 => (x"51",x"c1",x"c2",x"81"),
  1530 => (x"49",x"66",x"e8",x"c0"),
  1531 => (x"66",x"c4",x"81",x"c2"),
  1532 => (x"51",x"c0",x"81",x"bf"),
  1533 => (x"d0",x"c1",x"48",x"6e"),
  1534 => (x"49",x"6e",x"78",x"ce"),
  1535 => (x"66",x"d0",x"81",x"c8"),
  1536 => (x"c9",x"49",x"6e",x"51"),
  1537 => (x"51",x"66",x"d4",x"81"),
  1538 => (x"81",x"ca",x"49",x"6e"),
  1539 => (x"d0",x"51",x"66",x"dc"),
  1540 => (x"80",x"c1",x"48",x"66"),
  1541 => (x"48",x"58",x"a6",x"d4"),
  1542 => (x"78",x"c1",x"80",x"d8"),
  1543 => (x"ff",x"87",x"e8",x"c4"),
  1544 => (x"70",x"87",x"eb",x"dc"),
  1545 => (x"a6",x"ec",x"c0",x"49"),
  1546 => (x"e1",x"dc",x"ff",x"59"),
  1547 => (x"c0",x"49",x"70",x"87"),
  1548 => (x"dc",x"59",x"a6",x"e0"),
  1549 => (x"ec",x"c0",x"48",x"66"),
  1550 => (x"ca",x"c0",x"05",x"a8"),
  1551 => (x"48",x"a6",x"dc",x"87"),
  1552 => (x"78",x"66",x"e8",x"c0"),
  1553 => (x"ff",x"87",x"c4",x"c0"),
  1554 => (x"c8",x"87",x"d0",x"d9"),
  1555 => (x"91",x"cb",x"49",x"66"),
  1556 => (x"48",x"66",x"c0",x"c1"),
  1557 => (x"7e",x"70",x"80",x"71"),
  1558 => (x"82",x"c8",x"4a",x"6e"),
  1559 => (x"81",x"ca",x"49",x"6e"),
  1560 => (x"51",x"66",x"e8",x"c0"),
  1561 => (x"c1",x"49",x"66",x"dc"),
  1562 => (x"66",x"e8",x"c0",x"81"),
  1563 => (x"71",x"48",x"c1",x"89"),
  1564 => (x"c1",x"49",x"70",x"30"),
  1565 => (x"7a",x"97",x"71",x"89"),
  1566 => (x"bf",x"c0",x"f7",x"c2"),
  1567 => (x"66",x"e8",x"c0",x"49"),
  1568 => (x"4a",x"6a",x"97",x"29"),
  1569 => (x"c0",x"98",x"71",x"48"),
  1570 => (x"6e",x"58",x"a6",x"f0"),
  1571 => (x"69",x"81",x"c4",x"49"),
  1572 => (x"66",x"e0",x"c0",x"4d"),
  1573 => (x"a8",x"66",x"c4",x"48"),
  1574 => (x"87",x"c8",x"c0",x"02"),
  1575 => (x"c0",x"48",x"a6",x"c4"),
  1576 => (x"87",x"c5",x"c0",x"78"),
  1577 => (x"c1",x"48",x"a6",x"c4"),
  1578 => (x"1e",x"66",x"c4",x"78"),
  1579 => (x"75",x"1e",x"e0",x"c0"),
  1580 => (x"ea",x"d8",x"ff",x"49"),
  1581 => (x"70",x"86",x"c8",x"87"),
  1582 => (x"ac",x"b7",x"c0",x"4c"),
  1583 => (x"87",x"d4",x"c1",x"06"),
  1584 => (x"e0",x"c0",x"85",x"74"),
  1585 => (x"75",x"89",x"74",x"49"),
  1586 => (x"de",x"e7",x"c1",x"4b"),
  1587 => (x"df",x"fe",x"71",x"4a"),
  1588 => (x"85",x"c2",x"87",x"d6"),
  1589 => (x"48",x"66",x"e4",x"c0"),
  1590 => (x"e8",x"c0",x"80",x"c1"),
  1591 => (x"ec",x"c0",x"58",x"a6"),
  1592 => (x"81",x"c1",x"49",x"66"),
  1593 => (x"c0",x"02",x"a9",x"70"),
  1594 => (x"a6",x"c4",x"87",x"c8"),
  1595 => (x"c0",x"78",x"c0",x"48"),
  1596 => (x"a6",x"c4",x"87",x"c5"),
  1597 => (x"c4",x"78",x"c1",x"48"),
  1598 => (x"a4",x"c2",x"1e",x"66"),
  1599 => (x"48",x"e0",x"c0",x"49"),
  1600 => (x"49",x"70",x"88",x"71"),
  1601 => (x"ff",x"49",x"75",x"1e"),
  1602 => (x"c8",x"87",x"d4",x"d7"),
  1603 => (x"a8",x"b7",x"c0",x"86"),
  1604 => (x"87",x"c0",x"ff",x"01"),
  1605 => (x"02",x"66",x"e4",x"c0"),
  1606 => (x"6e",x"87",x"d1",x"c0"),
  1607 => (x"c0",x"81",x"c9",x"49"),
  1608 => (x"6e",x"51",x"66",x"e4"),
  1609 => (x"df",x"d2",x"c1",x"48"),
  1610 => (x"87",x"cc",x"c0",x"78"),
  1611 => (x"81",x"c9",x"49",x"6e"),
  1612 => (x"48",x"6e",x"51",x"c2"),
  1613 => (x"78",x"d3",x"d3",x"c1"),
  1614 => (x"48",x"a6",x"e8",x"c0"),
  1615 => (x"c6",x"c0",x"78",x"c1"),
  1616 => (x"c6",x"d6",x"ff",x"87"),
  1617 => (x"c0",x"4c",x"70",x"87"),
  1618 => (x"c0",x"02",x"66",x"e8"),
  1619 => (x"66",x"c8",x"87",x"f5"),
  1620 => (x"a8",x"66",x"cc",x"48"),
  1621 => (x"87",x"cb",x"c0",x"04"),
  1622 => (x"c1",x"48",x"66",x"c8"),
  1623 => (x"58",x"a6",x"cc",x"80"),
  1624 => (x"cc",x"87",x"e0",x"c0"),
  1625 => (x"88",x"c1",x"48",x"66"),
  1626 => (x"c0",x"58",x"a6",x"d0"),
  1627 => (x"c6",x"c1",x"87",x"d5"),
  1628 => (x"c8",x"c0",x"05",x"ac"),
  1629 => (x"48",x"66",x"d0",x"87"),
  1630 => (x"a6",x"d4",x"80",x"c1"),
  1631 => (x"ca",x"d5",x"ff",x"58"),
  1632 => (x"d4",x"4c",x"70",x"87"),
  1633 => (x"80",x"c1",x"48",x"66"),
  1634 => (x"74",x"58",x"a6",x"d8"),
  1635 => (x"cb",x"c0",x"02",x"9c"),
  1636 => (x"48",x"66",x"c8",x"87"),
  1637 => (x"a8",x"66",x"c8",x"c1"),
  1638 => (x"87",x"ef",x"f2",x"04"),
  1639 => (x"87",x"e2",x"d4",x"ff"),
  1640 => (x"c7",x"48",x"66",x"c8"),
  1641 => (x"e5",x"c0",x"03",x"a8"),
  1642 => (x"d4",x"f3",x"c2",x"87"),
  1643 => (x"c8",x"78",x"c0",x"48"),
  1644 => (x"91",x"cb",x"49",x"66"),
  1645 => (x"81",x"66",x"c0",x"c1"),
  1646 => (x"6a",x"4a",x"a1",x"c4"),
  1647 => (x"79",x"52",x"c0",x"4a"),
  1648 => (x"c1",x"48",x"66",x"c8"),
  1649 => (x"58",x"a6",x"cc",x"80"),
  1650 => (x"ff",x"04",x"a8",x"c7"),
  1651 => (x"d0",x"ff",x"87",x"db"),
  1652 => (x"f7",x"de",x"ff",x"8e"),
  1653 => (x"61",x"6f",x"4c",x"87"),
  1654 => (x"2e",x"2a",x"20",x"64"),
  1655 => (x"20",x"3a",x"00",x"20"),
  1656 => (x"1e",x"73",x"1e",x"00"),
  1657 => (x"02",x"9b",x"4b",x"71"),
  1658 => (x"f3",x"c2",x"87",x"c6"),
  1659 => (x"78",x"c0",x"48",x"d0"),
  1660 => (x"f3",x"c2",x"1e",x"c7"),
  1661 => (x"1e",x"49",x"bf",x"d0"),
  1662 => (x"1e",x"fd",x"ea",x"c1"),
  1663 => (x"bf",x"c4",x"f2",x"c2"),
  1664 => (x"87",x"ef",x"ed",x"49"),
  1665 => (x"f2",x"c2",x"86",x"cc"),
  1666 => (x"e9",x"49",x"bf",x"c4"),
  1667 => (x"9b",x"73",x"87",x"e9"),
  1668 => (x"c1",x"87",x"c8",x"02"),
  1669 => (x"c0",x"49",x"fd",x"ea"),
  1670 => (x"ff",x"87",x"c5",x"e4"),
  1671 => (x"1e",x"87",x"f1",x"dd"),
  1672 => (x"c1",x"87",x"d4",x"c7"),
  1673 => (x"87",x"f9",x"fe",x"49"),
  1674 => (x"87",x"c9",x"e4",x"fe"),
  1675 => (x"cd",x"02",x"98",x"70"),
  1676 => (x"c4",x"ed",x"fe",x"87"),
  1677 => (x"02",x"98",x"70",x"87"),
  1678 => (x"4a",x"c1",x"87",x"c4"),
  1679 => (x"4a",x"c0",x"87",x"c2"),
  1680 => (x"ce",x"05",x"9a",x"72"),
  1681 => (x"c1",x"1e",x"c0",x"87"),
  1682 => (x"c0",x"49",x"f0",x"e9"),
  1683 => (x"c4",x"87",x"d7",x"f0"),
  1684 => (x"c0",x"87",x"fe",x"86"),
  1685 => (x"fb",x"e9",x"c1",x"1e"),
  1686 => (x"c9",x"f0",x"c0",x"49"),
  1687 => (x"c0",x"1e",x"c0",x"87"),
  1688 => (x"70",x"87",x"cd",x"fa"),
  1689 => (x"fd",x"ef",x"c0",x"49"),
  1690 => (x"87",x"ca",x"c3",x"87"),
  1691 => (x"4f",x"26",x"8e",x"f8"),
  1692 => (x"66",x"20",x"44",x"53"),
  1693 => (x"65",x"6c",x"69",x"61"),
  1694 => (x"42",x"00",x"2e",x"64"),
  1695 => (x"69",x"74",x"6f",x"6f"),
  1696 => (x"2e",x"2e",x"67",x"6e"),
  1697 => (x"c0",x"1e",x"00",x"2e"),
  1698 => (x"c0",x"87",x"f1",x"e6"),
  1699 => (x"f6",x"87",x"de",x"f3"),
  1700 => (x"1e",x"4f",x"26",x"87"),
  1701 => (x"48",x"d0",x"f3",x"c2"),
  1702 => (x"f2",x"c2",x"78",x"c0"),
  1703 => (x"78",x"c0",x"48",x"c4"),
  1704 => (x"e1",x"87",x"fc",x"fd"),
  1705 => (x"26",x"48",x"c0",x"87"),
  1706 => (x"01",x"00",x"00",x"4f"),
  1707 => (x"80",x"00",x"00",x"00"),
  1708 => (x"69",x"78",x"45",x"20"),
  1709 => (x"20",x"80",x"00",x"74"),
  1710 => (x"6b",x"63",x"61",x"42"),
  1711 => (x"00",x"12",x"13",x"00"),
  1712 => (x"00",x"2c",x"e4",x"00"),
  1713 => (x"00",x"00",x"00",x"00"),
  1714 => (x"00",x"00",x"12",x"13"),
  1715 => (x"00",x"00",x"2d",x"02"),
  1716 => (x"13",x"00",x"00",x"00"),
  1717 => (x"20",x"00",x"00",x"12"),
  1718 => (x"00",x"00",x"00",x"2d"),
  1719 => (x"12",x"13",x"00",x"00"),
  1720 => (x"2d",x"3e",x"00",x"00"),
  1721 => (x"00",x"00",x"00",x"00"),
  1722 => (x"00",x"12",x"13",x"00"),
  1723 => (x"00",x"2d",x"5c",x"00"),
  1724 => (x"00",x"00",x"00",x"00"),
  1725 => (x"00",x"00",x"12",x"13"),
  1726 => (x"00",x"00",x"2d",x"7a"),
  1727 => (x"13",x"00",x"00",x"00"),
  1728 => (x"98",x"00",x"00",x"12"),
  1729 => (x"00",x"00",x"00",x"2d"),
  1730 => (x"14",x"4f",x"00",x"00"),
  1731 => (x"00",x"00",x"00",x"00"),
  1732 => (x"00",x"00",x"00",x"00"),
  1733 => (x"00",x"14",x"e4",x"00"),
  1734 => (x"00",x"00",x"00",x"00"),
  1735 => (x"00",x"00",x"00",x"00"),
  1736 => (x"48",x"f0",x"fe",x"1e"),
  1737 => (x"09",x"cd",x"78",x"c0"),
  1738 => (x"4f",x"26",x"09",x"79"),
  1739 => (x"f0",x"fe",x"1e",x"1e"),
  1740 => (x"26",x"48",x"7e",x"bf"),
  1741 => (x"fe",x"1e",x"4f",x"26"),
  1742 => (x"78",x"c1",x"48",x"f0"),
  1743 => (x"fe",x"1e",x"4f",x"26"),
  1744 => (x"78",x"c0",x"48",x"f0"),
  1745 => (x"71",x"1e",x"4f",x"26"),
  1746 => (x"52",x"52",x"c0",x"4a"),
  1747 => (x"5e",x"0e",x"4f",x"26"),
  1748 => (x"0e",x"5d",x"5c",x"5b"),
  1749 => (x"4d",x"71",x"86",x"f4"),
  1750 => (x"c1",x"7e",x"6d",x"97"),
  1751 => (x"6c",x"97",x"4c",x"a5"),
  1752 => (x"58",x"a6",x"c8",x"48"),
  1753 => (x"66",x"c4",x"48",x"6e"),
  1754 => (x"87",x"c5",x"05",x"a8"),
  1755 => (x"e6",x"c0",x"48",x"ff"),
  1756 => (x"87",x"ca",x"ff",x"87"),
  1757 => (x"97",x"49",x"a5",x"c2"),
  1758 => (x"a3",x"71",x"4b",x"6c"),
  1759 => (x"4b",x"6b",x"97",x"4b"),
  1760 => (x"6e",x"7e",x"6c",x"97"),
  1761 => (x"c8",x"80",x"c1",x"48"),
  1762 => (x"98",x"c7",x"58",x"a6"),
  1763 => (x"70",x"58",x"a6",x"cc"),
  1764 => (x"e1",x"fe",x"7c",x"97"),
  1765 => (x"f4",x"48",x"73",x"87"),
  1766 => (x"26",x"4d",x"26",x"8e"),
  1767 => (x"26",x"4b",x"26",x"4c"),
  1768 => (x"5b",x"5e",x"0e",x"4f"),
  1769 => (x"86",x"f4",x"0e",x"5c"),
  1770 => (x"66",x"d8",x"4c",x"71"),
  1771 => (x"9a",x"ff",x"c3",x"4a"),
  1772 => (x"97",x"4b",x"a4",x"c2"),
  1773 => (x"a1",x"73",x"49",x"6c"),
  1774 => (x"97",x"51",x"72",x"49"),
  1775 => (x"48",x"6e",x"7e",x"6c"),
  1776 => (x"a6",x"c8",x"80",x"c1"),
  1777 => (x"cc",x"98",x"c7",x"58"),
  1778 => (x"54",x"70",x"58",x"a6"),
  1779 => (x"ca",x"ff",x"8e",x"f4"),
  1780 => (x"fd",x"1e",x"1e",x"87"),
  1781 => (x"bf",x"e0",x"87",x"e8"),
  1782 => (x"e0",x"c0",x"49",x"4a"),
  1783 => (x"cb",x"02",x"99",x"c0"),
  1784 => (x"c2",x"1e",x"72",x"87"),
  1785 => (x"fe",x"49",x"f6",x"f6"),
  1786 => (x"86",x"c4",x"87",x"f7"),
  1787 => (x"70",x"87",x"fd",x"fc"),
  1788 => (x"87",x"c2",x"fd",x"7e"),
  1789 => (x"1e",x"4f",x"26",x"26"),
  1790 => (x"49",x"f6",x"f6",x"c2"),
  1791 => (x"c1",x"87",x"c7",x"fd"),
  1792 => (x"fc",x"49",x"d1",x"ef"),
  1793 => (x"f7",x"c3",x"87",x"da"),
  1794 => (x"0e",x"4f",x"26",x"87"),
  1795 => (x"5d",x"5c",x"5b",x"5e"),
  1796 => (x"c2",x"4d",x"71",x"0e"),
  1797 => (x"fc",x"49",x"f6",x"f6"),
  1798 => (x"4b",x"70",x"87",x"f4"),
  1799 => (x"04",x"ab",x"b7",x"c0"),
  1800 => (x"c3",x"87",x"c2",x"c3"),
  1801 => (x"c9",x"05",x"ab",x"f0"),
  1802 => (x"ef",x"f3",x"c1",x"87"),
  1803 => (x"c2",x"78",x"c1",x"48"),
  1804 => (x"e0",x"c3",x"87",x"e3"),
  1805 => (x"87",x"c9",x"05",x"ab"),
  1806 => (x"48",x"f3",x"f3",x"c1"),
  1807 => (x"d4",x"c2",x"78",x"c1"),
  1808 => (x"f3",x"f3",x"c1",x"87"),
  1809 => (x"87",x"c6",x"02",x"bf"),
  1810 => (x"4c",x"a3",x"c0",x"c2"),
  1811 => (x"4c",x"73",x"87",x"c2"),
  1812 => (x"bf",x"ef",x"f3",x"c1"),
  1813 => (x"87",x"e0",x"c0",x"02"),
  1814 => (x"b7",x"c4",x"49",x"74"),
  1815 => (x"f5",x"c1",x"91",x"29"),
  1816 => (x"4a",x"74",x"81",x"cf"),
  1817 => (x"92",x"c2",x"9a",x"cf"),
  1818 => (x"30",x"72",x"48",x"c1"),
  1819 => (x"ba",x"ff",x"4a",x"70"),
  1820 => (x"98",x"69",x"48",x"72"),
  1821 => (x"87",x"db",x"79",x"70"),
  1822 => (x"b7",x"c4",x"49",x"74"),
  1823 => (x"f5",x"c1",x"91",x"29"),
  1824 => (x"4a",x"74",x"81",x"cf"),
  1825 => (x"92",x"c2",x"9a",x"cf"),
  1826 => (x"30",x"72",x"48",x"c3"),
  1827 => (x"69",x"48",x"4a",x"70"),
  1828 => (x"75",x"79",x"70",x"b0"),
  1829 => (x"f0",x"c0",x"05",x"9d"),
  1830 => (x"48",x"d0",x"ff",x"87"),
  1831 => (x"ff",x"78",x"e1",x"c8"),
  1832 => (x"78",x"c5",x"48",x"d4"),
  1833 => (x"bf",x"f3",x"f3",x"c1"),
  1834 => (x"c3",x"87",x"c3",x"02"),
  1835 => (x"f3",x"c1",x"78",x"e0"),
  1836 => (x"c6",x"02",x"bf",x"ef"),
  1837 => (x"48",x"d4",x"ff",x"87"),
  1838 => (x"ff",x"78",x"f0",x"c3"),
  1839 => (x"78",x"73",x"48",x"d4"),
  1840 => (x"c8",x"48",x"d0",x"ff"),
  1841 => (x"e0",x"c0",x"78",x"e1"),
  1842 => (x"f3",x"f3",x"c1",x"78"),
  1843 => (x"c1",x"78",x"c0",x"48"),
  1844 => (x"c0",x"48",x"ef",x"f3"),
  1845 => (x"f6",x"f6",x"c2",x"78"),
  1846 => (x"87",x"f2",x"f9",x"49"),
  1847 => (x"b7",x"c0",x"4b",x"70"),
  1848 => (x"fe",x"fc",x"03",x"ab"),
  1849 => (x"26",x"48",x"c0",x"87"),
  1850 => (x"26",x"4c",x"26",x"4d"),
  1851 => (x"00",x"4f",x"26",x"4b"),
  1852 => (x"00",x"00",x"00",x"00"),
  1853 => (x"1e",x"00",x"00",x"00"),
  1854 => (x"fc",x"49",x"4a",x"71"),
  1855 => (x"4f",x"26",x"87",x"cd"),
  1856 => (x"72",x"4a",x"c0",x"1e"),
  1857 => (x"c1",x"91",x"c4",x"49"),
  1858 => (x"c0",x"81",x"cf",x"f5"),
  1859 => (x"d0",x"82",x"c1",x"79"),
  1860 => (x"ee",x"04",x"aa",x"b7"),
  1861 => (x"0e",x"4f",x"26",x"87"),
  1862 => (x"5d",x"5c",x"5b",x"5e"),
  1863 => (x"f8",x"4d",x"71",x"0e"),
  1864 => (x"4a",x"75",x"87",x"dc"),
  1865 => (x"92",x"2a",x"b7",x"c4"),
  1866 => (x"82",x"cf",x"f5",x"c1"),
  1867 => (x"9c",x"cf",x"4c",x"75"),
  1868 => (x"49",x"6a",x"94",x"c2"),
  1869 => (x"c3",x"2b",x"74",x"4b"),
  1870 => (x"74",x"48",x"c2",x"9b"),
  1871 => (x"ff",x"4c",x"70",x"30"),
  1872 => (x"71",x"48",x"74",x"bc"),
  1873 => (x"f7",x"7a",x"70",x"98"),
  1874 => (x"48",x"73",x"87",x"ec"),
  1875 => (x"00",x"87",x"d8",x"fe"),
  1876 => (x"00",x"00",x"00",x"00"),
  1877 => (x"00",x"00",x"00",x"00"),
  1878 => (x"00",x"00",x"00",x"00"),
  1879 => (x"00",x"00",x"00",x"00"),
  1880 => (x"00",x"00",x"00",x"00"),
  1881 => (x"00",x"00",x"00",x"00"),
  1882 => (x"00",x"00",x"00",x"00"),
  1883 => (x"00",x"00",x"00",x"00"),
  1884 => (x"00",x"00",x"00",x"00"),
  1885 => (x"00",x"00",x"00",x"00"),
  1886 => (x"00",x"00",x"00",x"00"),
  1887 => (x"00",x"00",x"00",x"00"),
  1888 => (x"00",x"00",x"00",x"00"),
  1889 => (x"00",x"00",x"00",x"00"),
  1890 => (x"00",x"00",x"00",x"00"),
  1891 => (x"1e",x"00",x"00",x"00"),
  1892 => (x"c8",x"48",x"d0",x"ff"),
  1893 => (x"48",x"71",x"78",x"e1"),
  1894 => (x"78",x"08",x"d4",x"ff"),
  1895 => (x"ff",x"1e",x"4f",x"26"),
  1896 => (x"e1",x"c8",x"48",x"d0"),
  1897 => (x"ff",x"48",x"71",x"78"),
  1898 => (x"c4",x"78",x"08",x"d4"),
  1899 => (x"d4",x"ff",x"48",x"66"),
  1900 => (x"4f",x"26",x"78",x"08"),
  1901 => (x"c4",x"4a",x"71",x"1e"),
  1902 => (x"72",x"1e",x"49",x"66"),
  1903 => (x"87",x"de",x"ff",x"49"),
  1904 => (x"c0",x"48",x"d0",x"ff"),
  1905 => (x"26",x"26",x"78",x"e0"),
  1906 => (x"1e",x"73",x"1e",x"4f"),
  1907 => (x"66",x"c8",x"4b",x"71"),
  1908 => (x"4a",x"73",x"1e",x"49"),
  1909 => (x"49",x"a2",x"e0",x"c1"),
  1910 => (x"26",x"87",x"d9",x"ff"),
  1911 => (x"4d",x"26",x"87",x"c4"),
  1912 => (x"4b",x"26",x"4c",x"26"),
  1913 => (x"73",x"1e",x"4f",x"26"),
  1914 => (x"4b",x"4a",x"71",x"1e"),
  1915 => (x"03",x"ab",x"b7",x"c2"),
  1916 => (x"49",x"a3",x"87",x"c8"),
  1917 => (x"9a",x"ff",x"c3",x"4a"),
  1918 => (x"a3",x"ce",x"87",x"c7"),
  1919 => (x"ff",x"c3",x"4a",x"49"),
  1920 => (x"49",x"66",x"c8",x"9a"),
  1921 => (x"fe",x"49",x"72",x"1e"),
  1922 => (x"ff",x"26",x"87",x"ea"),
  1923 => (x"ff",x"1e",x"87",x"d4"),
  1924 => (x"ff",x"c3",x"4a",x"d4"),
  1925 => (x"48",x"d0",x"ff",x"7a"),
  1926 => (x"de",x"78",x"e1",x"c0"),
  1927 => (x"c0",x"f7",x"c2",x"7a"),
  1928 => (x"48",x"49",x"7a",x"bf"),
  1929 => (x"7a",x"70",x"28",x"c8"),
  1930 => (x"28",x"d0",x"48",x"71"),
  1931 => (x"48",x"71",x"7a",x"70"),
  1932 => (x"7a",x"70",x"28",x"d8"),
  1933 => (x"c0",x"48",x"d0",x"ff"),
  1934 => (x"4f",x"26",x"78",x"e0"),
  1935 => (x"5c",x"5b",x"5e",x"0e"),
  1936 => (x"4c",x"71",x"0e",x"5d"),
  1937 => (x"bf",x"c0",x"f7",x"c2"),
  1938 => (x"29",x"74",x"49",x"4d"),
  1939 => (x"66",x"d0",x"4b",x"71"),
  1940 => (x"d4",x"83",x"c1",x"9b"),
  1941 => (x"04",x"ab",x"b7",x"66"),
  1942 => (x"4b",x"c0",x"87",x"c2"),
  1943 => (x"74",x"49",x"66",x"d0"),
  1944 => (x"75",x"b9",x"ff",x"31"),
  1945 => (x"74",x"4a",x"73",x"99"),
  1946 => (x"71",x"48",x"72",x"32"),
  1947 => (x"c4",x"f7",x"c2",x"b0"),
  1948 => (x"87",x"da",x"fe",x"58"),
  1949 => (x"4c",x"26",x"4d",x"26"),
  1950 => (x"4f",x"26",x"4b",x"26"),
  1951 => (x"48",x"d0",x"ff",x"1e"),
  1952 => (x"71",x"78",x"c9",x"c8"),
  1953 => (x"08",x"d4",x"ff",x"48"),
  1954 => (x"1e",x"4f",x"26",x"78"),
  1955 => (x"eb",x"49",x"4a",x"71"),
  1956 => (x"48",x"d0",x"ff",x"87"),
  1957 => (x"4f",x"26",x"78",x"c8"),
  1958 => (x"71",x"1e",x"73",x"1e"),
  1959 => (x"d0",x"f7",x"c2",x"4b"),
  1960 => (x"87",x"c3",x"02",x"bf"),
  1961 => (x"ff",x"87",x"eb",x"c2"),
  1962 => (x"c9",x"c8",x"48",x"d0"),
  1963 => (x"c0",x"49",x"73",x"78"),
  1964 => (x"d4",x"ff",x"b1",x"e0"),
  1965 => (x"c2",x"78",x"71",x"48"),
  1966 => (x"c0",x"48",x"c4",x"f7"),
  1967 => (x"02",x"66",x"c8",x"78"),
  1968 => (x"ff",x"c3",x"87",x"c5"),
  1969 => (x"c0",x"87",x"c2",x"49"),
  1970 => (x"cc",x"f7",x"c2",x"49"),
  1971 => (x"02",x"66",x"cc",x"59"),
  1972 => (x"d5",x"c5",x"87",x"c6"),
  1973 => (x"87",x"c4",x"4a",x"d5"),
  1974 => (x"4a",x"ff",x"ff",x"cf"),
  1975 => (x"5a",x"d0",x"f7",x"c2"),
  1976 => (x"48",x"d0",x"f7",x"c2"),
  1977 => (x"87",x"c4",x"78",x"c1"),
  1978 => (x"4c",x"26",x"4d",x"26"),
  1979 => (x"4f",x"26",x"4b",x"26"),
  1980 => (x"5c",x"5b",x"5e",x"0e"),
  1981 => (x"4a",x"71",x"0e",x"5d"),
  1982 => (x"bf",x"cc",x"f7",x"c2"),
  1983 => (x"02",x"9a",x"72",x"4c"),
  1984 => (x"c8",x"49",x"87",x"cb"),
  1985 => (x"ce",x"fa",x"c1",x"91"),
  1986 => (x"c4",x"83",x"71",x"4b"),
  1987 => (x"ce",x"fe",x"c1",x"87"),
  1988 => (x"13",x"4d",x"c0",x"4b"),
  1989 => (x"c2",x"99",x"74",x"49"),
  1990 => (x"b9",x"bf",x"c8",x"f7"),
  1991 => (x"71",x"48",x"d4",x"ff"),
  1992 => (x"2c",x"b7",x"c1",x"78"),
  1993 => (x"ad",x"b7",x"c8",x"85"),
  1994 => (x"c2",x"87",x"e8",x"04"),
  1995 => (x"48",x"bf",x"c4",x"f7"),
  1996 => (x"f7",x"c2",x"80",x"c8"),
  1997 => (x"ef",x"fe",x"58",x"c8"),
  1998 => (x"1e",x"73",x"1e",x"87"),
  1999 => (x"4a",x"13",x"4b",x"71"),
  2000 => (x"87",x"cb",x"02",x"9a"),
  2001 => (x"e7",x"fe",x"49",x"72"),
  2002 => (x"9a",x"4a",x"13",x"87"),
  2003 => (x"fe",x"87",x"f5",x"05"),
  2004 => (x"c2",x"1e",x"87",x"da"),
  2005 => (x"49",x"bf",x"c4",x"f7"),
  2006 => (x"48",x"c4",x"f7",x"c2"),
  2007 => (x"c4",x"78",x"a1",x"c1"),
  2008 => (x"03",x"a9",x"b7",x"c0"),
  2009 => (x"d4",x"ff",x"87",x"db"),
  2010 => (x"c8",x"f7",x"c2",x"48"),
  2011 => (x"f7",x"c2",x"78",x"bf"),
  2012 => (x"c2",x"49",x"bf",x"c4"),
  2013 => (x"c1",x"48",x"c4",x"f7"),
  2014 => (x"c0",x"c4",x"78",x"a1"),
  2015 => (x"e5",x"04",x"a9",x"b7"),
  2016 => (x"48",x"d0",x"ff",x"87"),
  2017 => (x"f7",x"c2",x"78",x"c8"),
  2018 => (x"78",x"c0",x"48",x"d0"),
  2019 => (x"00",x"00",x"4f",x"26"),
  2020 => (x"00",x"00",x"00",x"00"),
  2021 => (x"00",x"00",x"00",x"00"),
  2022 => (x"00",x"5f",x"5f",x"00"),
  2023 => (x"03",x"00",x"00",x"00"),
  2024 => (x"03",x"03",x"00",x"03"),
  2025 => (x"7f",x"14",x"00",x"00"),
  2026 => (x"7f",x"7f",x"14",x"7f"),
  2027 => (x"24",x"00",x"00",x"14"),
  2028 => (x"3a",x"6b",x"6b",x"2e"),
  2029 => (x"6a",x"4c",x"00",x"12"),
  2030 => (x"56",x"6c",x"18",x"36"),
  2031 => (x"7e",x"30",x"00",x"32"),
  2032 => (x"3a",x"77",x"59",x"4f"),
  2033 => (x"00",x"00",x"40",x"68"),
  2034 => (x"00",x"03",x"07",x"04"),
  2035 => (x"00",x"00",x"00",x"00"),
  2036 => (x"41",x"63",x"3e",x"1c"),
  2037 => (x"00",x"00",x"00",x"00"),
  2038 => (x"1c",x"3e",x"63",x"41"),
  2039 => (x"2a",x"08",x"00",x"00"),
  2040 => (x"3e",x"1c",x"1c",x"3e"),
  2041 => (x"08",x"00",x"08",x"2a"),
  2042 => (x"08",x"3e",x"3e",x"08"),
  2043 => (x"00",x"00",x"00",x"08"),
  2044 => (x"00",x"60",x"e0",x"80"),
  2045 => (x"08",x"00",x"00",x"00"),
  2046 => (x"08",x"08",x"08",x"08"),
  2047 => (x"00",x"00",x"00",x"08"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

