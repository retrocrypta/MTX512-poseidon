library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom2 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom2 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"00606000",
     1 => x"60400000",
     2 => x"060c1830",
     3 => x"3e000103",
     4 => x"7f4d597f",
     5 => x"0400003e",
     6 => x"007f7f06",
     7 => x"42000000",
     8 => x"4f597163",
     9 => x"22000046",
    10 => x"7f494963",
    11 => x"1c180036",
    12 => x"7f7f1316",
    13 => x"27000010",
    14 => x"7d454567",
    15 => x"3c000039",
    16 => x"79494b7e",
    17 => x"01000030",
    18 => x"0f797101",
    19 => x"36000007",
    20 => x"7f49497f",
    21 => x"06000036",
    22 => x"3f69494f",
    23 => x"0000001e",
    24 => x"00666600",
    25 => x"00000000",
    26 => x"0066e680",
    27 => x"08000000",
    28 => x"22141408",
    29 => x"14000022",
    30 => x"14141414",
    31 => x"22000014",
    32 => x"08141422",
    33 => x"02000008",
    34 => x"0f595103",
    35 => x"7f3e0006",
    36 => x"1f555d41",
    37 => x"7e00001e",
    38 => x"7f09097f",
    39 => x"7f00007e",
    40 => x"7f49497f",
    41 => x"1c000036",
    42 => x"4141633e",
    43 => x"7f000041",
    44 => x"3e63417f",
    45 => x"7f00001c",
    46 => x"4149497f",
    47 => x"7f000041",
    48 => x"0109097f",
    49 => x"3e000001",
    50 => x"7b49417f",
    51 => x"7f00007a",
    52 => x"7f08087f",
    53 => x"0000007f",
    54 => x"417f7f41",
    55 => x"20000000",
    56 => x"7f404060",
    57 => x"7f7f003f",
    58 => x"63361c08",
    59 => x"7f000041",
    60 => x"4040407f",
    61 => x"7f7f0040",
    62 => x"7f060c06",
    63 => x"7f7f007f",
    64 => x"7f180c06",
    65 => x"3e00007f",
    66 => x"7f41417f",
    67 => x"7f00003e",
    68 => x"0f09097f",
    69 => x"7f3e0006",
    70 => x"7e7f6141",
    71 => x"7f000040",
    72 => x"7f19097f",
    73 => x"26000066",
    74 => x"7b594d6f",
    75 => x"01000032",
    76 => x"017f7f01",
    77 => x"3f000001",
    78 => x"7f40407f",
    79 => x"0f00003f",
    80 => x"3f70703f",
    81 => x"7f7f000f",
    82 => x"7f301830",
    83 => x"6341007f",
    84 => x"361c1c36",
    85 => x"03014163",
    86 => x"067c7c06",
    87 => x"71610103",
    88 => x"43474d59",
    89 => x"00000041",
    90 => x"41417f7f",
    91 => x"03010000",
    92 => x"30180c06",
    93 => x"00004060",
    94 => x"7f7f4141",
    95 => x"0c080000",
    96 => x"0c060306",
    97 => x"80800008",
    98 => x"80808080",
    99 => x"00000080",
   100 => x"04070300",
   101 => x"20000000",
   102 => x"7c545474",
   103 => x"7f000078",
   104 => x"7c44447f",
   105 => x"38000038",
   106 => x"4444447c",
   107 => x"38000000",
   108 => x"7f44447c",
   109 => x"3800007f",
   110 => x"5c54547c",
   111 => x"04000018",
   112 => x"05057f7e",
   113 => x"18000000",
   114 => x"fca4a4bc",
   115 => x"7f00007c",
   116 => x"7c04047f",
   117 => x"00000078",
   118 => x"407d3d00",
   119 => x"80000000",
   120 => x"7dfd8080",
   121 => x"7f000000",
   122 => x"6c38107f",
   123 => x"00000044",
   124 => x"407f3f00",
   125 => x"7c7c0000",
   126 => x"7c0c180c",
   127 => x"7c000078",
   128 => x"7c04047c",
   129 => x"38000078",
   130 => x"7c44447c",
   131 => x"fc000038",
   132 => x"3c2424fc",
   133 => x"18000018",
   134 => x"fc24243c",
   135 => x"7c0000fc",
   136 => x"0c04047c",
   137 => x"48000008",
   138 => x"7454545c",
   139 => x"04000020",
   140 => x"44447f3f",
   141 => x"3c000000",
   142 => x"7c40407c",
   143 => x"1c00007c",
   144 => x"3c60603c",
   145 => x"7c3c001c",
   146 => x"7c603060",
   147 => x"6c44003c",
   148 => x"6c381038",
   149 => x"1c000044",
   150 => x"3c60e0bc",
   151 => x"4400001c",
   152 => x"4c5c7464",
   153 => x"08000044",
   154 => x"41773e08",
   155 => x"00000041",
   156 => x"007f7f00",
   157 => x"41000000",
   158 => x"083e7741",
   159 => x"01020008",
   160 => x"02020301",
   161 => x"7f7f0001",
   162 => x"7f7f7f7f",
   163 => x"0808007f",
   164 => x"3e3e1c1c",
   165 => x"7f7f7f7f",
   166 => x"1c1c3e3e",
   167 => x"10000808",
   168 => x"187c7c18",
   169 => x"10000010",
   170 => x"307c7c30",
   171 => x"30100010",
   172 => x"1e786060",
   173 => x"66420006",
   174 => x"663c183c",
   175 => x"38780042",
   176 => x"6cc6c26a",
   177 => x"00600038",
   178 => x"00006000",
   179 => x"5e0e0060",
   180 => x"0e5d5c5b",
   181 => x"c24c711e",
   182 => x"4dbfe1f7",
   183 => x"1ec04bc0",
   184 => x"c702ab74",
   185 => x"48a6c487",
   186 => x"87c578c0",
   187 => x"c148a6c4",
   188 => x"1e66c478",
   189 => x"dfee4973",
   190 => x"c086c887",
   191 => x"efef49e0",
   192 => x"4aa5c487",
   193 => x"f0f0496a",
   194 => x"87c6f187",
   195 => x"83c185cb",
   196 => x"04abb7c8",
   197 => x"2687c7ff",
   198 => x"4c264d26",
   199 => x"4f264b26",
   200 => x"c24a711e",
   201 => x"c25ae5f7",
   202 => x"c748e5f7",
   203 => x"ddfe4978",
   204 => x"1e4f2687",
   205 => x"4a711e73",
   206 => x"03aab7c0",
   207 => x"dbc287d3",
   208 => x"c405bfcc",
   209 => x"c24bc187",
   210 => x"c24bc087",
   211 => x"c45bd0db",
   212 => x"d0dbc287",
   213 => x"ccdbc25a",
   214 => x"9ac14abf",
   215 => x"49a2c0c1",
   216 => x"fc87e8ec",
   217 => x"ccdbc248",
   218 => x"effe78bf",
   219 => x"4a711e87",
   220 => x"721e66c4",
   221 => x"87eee949",
   222 => x"1e4f2626",
   223 => x"bfccdbc2",
   224 => x"87f3e549",
   225 => x"48d9f7c2",
   226 => x"c278bfe8",
   227 => x"ec48d5f7",
   228 => x"f7c278bf",
   229 => x"494abfd9",
   230 => x"c899ffc3",
   231 => x"48722ab7",
   232 => x"f7c2b071",
   233 => x"4f2658e1",
   234 => x"5c5b5e0e",
   235 => x"4b710e5d",
   236 => x"c287c8ff",
   237 => x"c048d4f7",
   238 => x"e5497350",
   239 => x"497087d9",
   240 => x"cb9cc24c",
   241 => x"cbcc49ee",
   242 => x"4d497087",
   243 => x"97d4f7c2",
   244 => x"e2c105bf",
   245 => x"4966d087",
   246 => x"bfddf7c2",
   247 => x"87d60599",
   248 => x"c24966d4",
   249 => x"99bfd5f7",
   250 => x"7387cb05",
   251 => x"87e7e449",
   252 => x"c1029870",
   253 => x"4cc187c1",
   254 => x"7587c0fe",
   255 => x"87e0cb49",
   256 => x"c6029870",
   257 => x"d4f7c287",
   258 => x"c250c148",
   259 => x"bf97d4f7",
   260 => x"87e3c005",
   261 => x"bfddf7c2",
   262 => x"9966d049",
   263 => x"87d6ff05",
   264 => x"bfd5f7c2",
   265 => x"9966d449",
   266 => x"87caff05",
   267 => x"e6e34973",
   268 => x"05987087",
   269 => x"7487fffe",
   270 => x"87dcfb48",
   271 => x"5c5b5e0e",
   272 => x"86f40e5d",
   273 => x"ec4c4dc0",
   274 => x"a6c47ebf",
   275 => x"e1f7c248",
   276 => x"1ec178bf",
   277 => x"49c71ec0",
   278 => x"c887cdfd",
   279 => x"02987086",
   280 => x"49ff87cd",
   281 => x"c187ccfb",
   282 => x"eae249da",
   283 => x"c24dc187",
   284 => x"bf97d4f7",
   285 => x"d187c302",
   286 => x"f7c287c9",
   287 => x"c24bbfd9",
   288 => x"05bfccdb",
   289 => x"c487d9c1",
   290 => x"c0c848a6",
   291 => x"dac278c0",
   292 => x"976e7ef8",
   293 => x"486e49bf",
   294 => x"7e7080c1",
   295 => x"87f7e171",
   296 => x"c3029870",
   297 => x"b366c487",
   298 => x"c14866c4",
   299 => x"a6c828b7",
   300 => x"05987058",
   301 => x"c387dbff",
   302 => x"dae149fd",
   303 => x"49fac387",
   304 => x"7387d4e1",
   305 => x"99ffc349",
   306 => x"49c01e71",
   307 => x"7387defa",
   308 => x"29b7c849",
   309 => x"49c11e71",
   310 => x"c887d2fa",
   311 => x"87c1c686",
   312 => x"bfddf7c2",
   313 => x"dd029b4b",
   314 => x"c8dbc287",
   315 => x"efc749bf",
   316 => x"05987087",
   317 => x"4bc087c4",
   318 => x"e0c287d2",
   319 => x"87d4c749",
   320 => x"58ccdbc2",
   321 => x"dbc287c6",
   322 => x"78c048c8",
   323 => x"99c24973",
   324 => x"c387ce05",
   325 => x"dfff49eb",
   326 => x"497087fd",
   327 => x"c20299c2",
   328 => x"734cfb87",
   329 => x"0599c149",
   330 => x"f4c387ce",
   331 => x"e6dfff49",
   332 => x"c2497087",
   333 => x"87c20299",
   334 => x"49734cfa",
   335 => x"ce0599c8",
   336 => x"49f5c387",
   337 => x"87cfdfff",
   338 => x"99c24970",
   339 => x"c287d502",
   340 => x"02bfe5f7",
   341 => x"c14887ca",
   342 => x"e9f7c288",
   343 => x"87c2c058",
   344 => x"4dc14cff",
   345 => x"99c44973",
   346 => x"c387ce05",
   347 => x"deff49f2",
   348 => x"497087e5",
   349 => x"dc0299c2",
   350 => x"e5f7c287",
   351 => x"c7487ebf",
   352 => x"c003a8b7",
   353 => x"486e87cb",
   354 => x"f7c280c1",
   355 => x"c2c058e9",
   356 => x"c14cfe87",
   357 => x"49fdc34d",
   358 => x"87fbddff",
   359 => x"99c24970",
   360 => x"87d5c002",
   361 => x"bfe5f7c2",
   362 => x"87c9c002",
   363 => x"48e5f7c2",
   364 => x"c2c078c0",
   365 => x"c14cfd87",
   366 => x"49fac34d",
   367 => x"87d7ddff",
   368 => x"99c24970",
   369 => x"87d9c002",
   370 => x"bfe5f7c2",
   371 => x"a8b7c748",
   372 => x"87c9c003",
   373 => x"48e5f7c2",
   374 => x"c2c078c7",
   375 => x"c14cfc87",
   376 => x"acb7c04d",
   377 => x"87d1c003",
   378 => x"c14a66c4",
   379 => x"026a82d8",
   380 => x"6a87c6c0",
   381 => x"7349744b",
   382 => x"c31ec00f",
   383 => x"dac11ef0",
   384 => x"87e4f649",
   385 => x"987086c8",
   386 => x"87e2c002",
   387 => x"c248a6c8",
   388 => x"78bfe5f7",
   389 => x"cb4966c8",
   390 => x"4866c491",
   391 => x"7e708071",
   392 => x"c002bf6e",
   393 => x"bf6e87c8",
   394 => x"4966c84b",
   395 => x"9d750f73",
   396 => x"87c8c002",
   397 => x"bfe5f7c2",
   398 => x"87d2f249",
   399 => x"bfd0dbc2",
   400 => x"87ddc002",
   401 => x"87d8c249",
   402 => x"c0029870",
   403 => x"f7c287d3",
   404 => x"f149bfe5",
   405 => x"49c087f8",
   406 => x"c287d8f3",
   407 => x"c048d0db",
   408 => x"f28ef478",
   409 => x"5e0e87f2",
   410 => x"0e5d5c5b",
   411 => x"c24c711e",
   412 => x"49bfe1f7",
   413 => x"4da1cdc1",
   414 => x"6981d1c1",
   415 => x"029c747e",
   416 => x"a5c487cf",
   417 => x"c27b744b",
   418 => x"49bfe1f7",
   419 => x"6e87d1f2",
   420 => x"059c747b",
   421 => x"4bc087c4",
   422 => x"4bc187c2",
   423 => x"d2f24973",
   424 => x"0266d487",
   425 => x"c04987c8",
   426 => x"4a7087ea",
   427 => x"4ac087c2",
   428 => x"5ad4dbc2",
   429 => x"87e0f126",
   430 => x"14111258",
   431 => x"231c1b1d",
   432 => x"9491595a",
   433 => x"f4ebf2f5",
   434 => x"00000000",
   435 => x"00000000",
   436 => x"00000000",
   437 => x"ff4a711e",
   438 => x"7249bfc8",
   439 => x"4f2648a1",
   440 => x"bfc8ff1e",
   441 => x"c0c0fe89",
   442 => x"a9c0c0c0",
   443 => x"c087c401",
   444 => x"c187c24a",
   445 => x"2648724a",
   446 => x"5b5e0e4f",
   447 => x"710e5d5c",
   448 => x"4cd4ff4b",
   449 => x"c04866d0",
   450 => x"ff49d678",
   451 => x"c387c0da",
   452 => x"496c7cff",
   453 => x"7199ffc3",
   454 => x"f0c3494d",
   455 => x"a9e0c199",
   456 => x"c387cb05",
   457 => x"486c7cff",
   458 => x"66d098c3",
   459 => x"ffc37808",
   460 => x"494a6c7c",
   461 => x"ffc331c8",
   462 => x"714a6c7c",
   463 => x"c84972b2",
   464 => x"7cffc331",
   465 => x"b2714a6c",
   466 => x"31c84972",
   467 => x"6c7cffc3",
   468 => x"ffb2714a",
   469 => x"e0c048d0",
   470 => x"029b7378",
   471 => x"7b7287c2",
   472 => x"4d264875",
   473 => x"4b264c26",
   474 => x"261e4f26",
   475 => x"5b5e0e4f",
   476 => x"86f80e5c",
   477 => x"a6c81e76",
   478 => x"87fdfd49",
   479 => x"4b7086c4",
   480 => x"a8c4486e",
   481 => x"87f4c203",
   482 => x"f0c34a73",
   483 => x"aad0c19a",
   484 => x"c187c702",
   485 => x"c205aae0",
   486 => x"497387e2",
   487 => x"c30299c8",
   488 => x"87c6ff87",
   489 => x"9cc34c73",
   490 => x"c105acc2",
   491 => x"66c487c4",
   492 => x"7131c949",
   493 => x"4a66c41e",
   494 => x"c292c8c1",
   495 => x"7249e9f7",
   496 => x"d7cdfe81",
   497 => x"ff49d887",
   498 => x"c887c4d7",
   499 => x"e5c21ec0",
   500 => x"e5fd49d2",
   501 => x"d0ff87ee",
   502 => x"78e0c048",
   503 => x"1ed2e5c2",
   504 => x"c14a66cc",
   505 => x"f7c292c8",
   506 => x"817249e9",
   507 => x"87ecc8fe",
   508 => x"acc186cc",
   509 => x"87c4c105",
   510 => x"c94966c4",
   511 => x"c41e7131",
   512 => x"c8c14a66",
   513 => x"e9f7c292",
   514 => x"fe817249",
   515 => x"c287cdcc",
   516 => x"c81ed2e5",
   517 => x"c8c14a66",
   518 => x"e9f7c292",
   519 => x"fe817249",
   520 => x"d787eac6",
   521 => x"e6d5ff49",
   522 => x"1ec0c887",
   523 => x"49d2e5c2",
   524 => x"87e9e3fd",
   525 => x"d0ff86cc",
   526 => x"78e0c048",
   527 => x"e3fc8ef8",
   528 => x"5b5e0e87",
   529 => x"1e0e5d5c",
   530 => x"d4ff4d71",
   531 => x"7e66d44c",
   532 => x"a8b7c348",
   533 => x"c087c506",
   534 => x"87e3c148",
   535 => x"dcfe4975",
   536 => x"1e7587d5",
   537 => x"c14b66c4",
   538 => x"f7c293c8",
   539 => x"497383e9",
   540 => x"87f2fffd",
   541 => x"4b6b83c8",
   542 => x"c848d0ff",
   543 => x"7cdd78e1",
   544 => x"ffc34973",
   545 => x"737c7199",
   546 => x"29b7c849",
   547 => x"7199ffc3",
   548 => x"d049737c",
   549 => x"ffc329b7",
   550 => x"737c7199",
   551 => x"29b7d849",
   552 => x"7cc07c71",
   553 => x"7c7c7c7c",
   554 => x"7c7c7c7c",
   555 => x"c07c7c7c",
   556 => x"66c478e0",
   557 => x"ff49dc1e",
   558 => x"c887f9d3",
   559 => x"26487386",
   560 => x"1e87dffa",
   561 => x"bfece3c2",
   562 => x"c2b9c149",
   563 => x"ff59f0e3",
   564 => x"ffc348d4",
   565 => x"48d0ff78",
   566 => x"ff78e1c0",
   567 => x"78c148d4",
   568 => x"787131c4",
   569 => x"c048d0ff",
   570 => x"4f2678e0",
   571 => x"00000000",
   572 => x"c21ec01e",
   573 => x"49bfc9e4",
   574 => x"c287c6fd",
   575 => x"49bfcde4",
   576 => x"87d9ddfe",
   577 => x"262648c0",
   578 => x"0029114f",
   579 => x"00291d00",
   580 => x"58544d00",
   581 => x"20323135",
   582 => x"44485620",
   583 => x"58544d00",
   584 => x"20323135",
   585 => x"4d4f5220",
   586 => x"4d4f5200",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
